module CCGRCG187( x0, x1, x2, x3, x4, x5, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17, f18, f19 );

	input x0, x1, x2, x3, x4, x5;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17, f18, f19;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269;

	not (d1, x1);
	not (d2, x2);
	buf (d3, x4);
	not (d4, x3);
	nor (d5, x1);
	and (d6, x0);
	nand (d7, x3, x4);
	not (d8, x4);
	xnor (d9, x0, x2);
	nor (d10, x0, x4);
	nor (d11, x0, x1);
	or (d12, x2, x3);
	xor (d13, x3, x4);
	buf (d14, x3);
	and (d15, x1, x2);
	nand (d16, x1, x5);
	nand (d17, x0, x1);
	and (d18, x1, x3);
	xnor (d19, x3, x5);
	and (d20, x5);
	or (d21, x2);
	xnor (d22, x3);
	xnor (d23, x0, x5);
	or (d24, x3);
	buf (d25, x1);
	not (d26, x0);
	xnor (d27, x2, x3);
	xnor (d28, x4, x5);
	nand (d29, x1, x4);
	nand (d30, x0, x2);
	nor (d31, x1, x2);
	xor (d32, d2, d29);
	not (d33, d14);
	nor (d34, d13, d18);
	buf (d35, d19);
	buf (d36, d22);
	xor (d37, d21, d23);
	or (d38, d14, d26);
	and (d39, d4, d27);
	nor (d40, d3, d25);
	and (d41, d1, d13);
	or (d42, d1, d22);
	xor (d43, d2, d14);
	not (d44, d29);
	nand (d45, d21, d28);
	nor (d46, d3, d24);
	or (d47, d5, d19);
	not (d48, d23);
	and (d49, d4, d21);
	not (d50, d27);
	buf (d51, d14);
	xnor (d52, d13, d30);
	or (d53, d19, d29);
	nand (d54, d22, d28);
	nand (d55, d28, d31);
	nor (d56, d18, d31);
	nand (d57, d4, d21);
	xor (d58, d15, d24);
	not (d59, d31);
	and (d60, d6, d20);
	xnor (d61, d13, d21);
	not (d62, d8);
	buf (d63, d12);
	not (d64, d7);
	nand (d65, d1, d2);
	or (d66, d4, d29);
	and (d67, d9, d31);
	xnor (d68, d3, d26);
	nor (d69, d20, d31);
	xor (d70, d2, d13);
	buf (d71, x0);
	xor (d72, d35, d53);
	and (d73, d36, d56);
	xor (d74, d36, d53);
	xor (d75, d63, d64);
	xor (d76, d43, d45);
	and (d77, d39, d56);
	nand (d78, d52, d59);
	xnor (d79, d41, d69);
	buf (d80, d51);
	nor (d81, d36, d58);
	nor (d82, d39, d44);
	nand (d83, d49, d56);
	xnor (d84, d59, d60);
	and (d85, d43, d45);
	xnor (d86, d45, d53);
	nor (d87, d42, d60);
	buf (d88, d37);
	xor (d89, d61, d64);
	or (d90, d36, d60);
	or (d91, d45, d56);
	xor (d92, d76, d80);
	not (d93, d24);
	and (d94, d76, d78);
	nand (d95, d75, d77);
	or (d96, d73, d86);
	nor (d97, d78, d86);
	not (d98, d12);
	nand (d99, d73, d91);
	buf (d100, d44);
	nand (d101, d82, d83);
	or (d102, d79, d87);
	nor (d103, d85, d88);
	and (d104, d85, d86);
	or (d105, d73, d77);
	nor (d106, d74, d79);
	xor (d107, d72, d73);
	not (d108, d69);
	nand (d109, d76, d85);
	xor (d110, d76, d81);
	xnor (d111, d75, d91);
	xor (d112, d81, d91);
	xor (d113, d77, d91);
	and (d114, d75, d90);
	not (d115, d22);
	xnor (d116, d74, d89);
	nor (d117, d72, d84);
	nand (d118, d77, d81);
	nand (d119, d74, d76);
	xnor (d120, d74, d88);
	nor (d121, d77, d86);
	xnor (d122, d75, d88);
	and (d123, d79, d90);
	nand (d124, d77, d87);
	nand (d125, d84, d87);
	nand (d126, d81, d91);
	buf (d127, d75);
	or (d128, d88, d89);
	nand (d129, d79, d83);
	and (d130, d72, d83);
	xnor (d131, d79, d83);
	or (d132, d72, d80);
	and (d133, d75, d82);
	nor (d134, d74, d91);
	xnor (d135, d76, d79);
	nand (d136, d78, d87);
	and (d137, d82, d88);
	or (d138, d73, d89);
	or (d139, d73, d89);
	xnor (d140, d73, d74);
	and (d141, d73, d79);
	xnor (d142, d84, d87);
	nor (d143, d78, d81);
	not (d144, d51);
	nand (d145, d84, d90);
	nor (d146, d73, d85);
	xor (d147, d72, d74);
	xnor (d148, d72, d85);
	xor (d149, d73, d85);
	xor (d150, d82, d91);
	nor (d151, d84);
	nand (d152, d72, d88);
	xor (d153, d87, d88);
	nor (d154, d83, d89);
	nand (d155, d75, d82);
	nand (d156, d74);
	xor (d157, d84, d88);
	xnor (d158, d74, d78);
	not (d159, d9);
	xor (d160, d79, d82);
	not (d161, d85);
	xnor (d162, d81, d83);
	buf (d163, d21);
	nor (d164, d72, d73);
	xnor (d165, d76, d91);
	nand (d166, d83, d84);
	xor (d167, d76, d81);
	xor (d168, d75, d79);
	nor (d169, d85, d86);
	and (d170, d79, d86);
	xnor (d171, d74, d86);
	xor (d172, d76, d85);
	buf (d173, d57);
	not (d174, d20);
	xor (d175, d80, d82);
	not (d176, d65);
	not (d177, d60);
	buf (d178, d105);
	or (d179, d161, d167);
	xnor (d180, d160, d176);
	buf (d181, d113);
	xor (d182, d94, d172);
	and (d183, d96, d119);
	xor (d184, d156, d174);
	buf (d185, d42);
	xnor (d186, d153, d174);
	nand (d187, d98, d110);
	nor (d188, d108, d136);
	or (d189, d127, d147);
	buf (d190, d54);
	or (d191, d117, d166);
	xnor (d192, d165, d173);
	nand (d193, d143, d176);
	nand (d194, d130, d176);
	or (d195, d102, d147);
	nor (d196, d141, d159);
	buf (d197, d159);
	not (d198, d25);
	nand (d199, d135, d174);
	xnor (d200, d111, d140);
	nand (d201, d99, d152);
	or (d202, d149, d163);
	not (d203, d36);
	not (d204, d58);
	xor (d205, d98, d137);
	nor (d206, d134, d175);
	xnor (d207, d139, d176);
	nand (d208, d94, d144);
	and (d209, d105, d140);
	xor (d210, d96, d108);
	or (d211, d130, d137);
	nor (d212, d106, d127);
	or (d213, d138, d170);
	nor (d214, d92, d96);
	nand (d215, d111, d150);
	xor (d216, d128, d165);
	or (d217, d111, d142);
	not (d218, d16);
	xor (d219, d100, d132);
	or (d220, d117, d135);
	xor (d221, d116, d118);
	nor (d222, d159, d161);
	and (d223, d132, d169);
	nand (d224, d94, d144);
	nand (d225, d103, d123);
	and (d226, d93, d120);
	nand (d227, d103, d110);
	nor (d228, d137, d171);
	nor (d229, d97, d129);
	or (d230, d142, d171);
	xor (d231, d97, d101);
	and (d232, d131, d152);
	and (d233, d103, d104);
	or (d234, d93, d105);
	buf (d235, d114);
	or (d236, d94, d125);
	or (d237, d109, d129);
	xnor (d238, d115, d121);
	not (d239, d124);
	xnor (d240, d118);
	nand (d241, d120, d147);
	xnor (d242, d164, d174);
	nor (d243, d129, d145);
	xnor (d244, d121, d170);
	xor (d245, d112, d119);
	buf (d246, d77);
	nand (d247, d126, d163);
	and (d248, d137, d161);
	or (d249, d113, d127);
	xor (d250, d98, d135);
	xor (d251, d95, d124);
	xor (d252, d99, d136);
	and (d253, d95, d101);
	or (d254, d113, d120);
	or (d255, d113, d162);
	nor (d256, d121, d161);
	and (d257, d107, d171);
	nand (d258, d145, d160);
	or (d259, d103, d164);
	or (d260, d100, d149);
	xor (d261, d110, d116);
	or (d262, d108, d140);
	xnor (d263, d117, d164);
	not (d264, d103);
	nand (d265, d164, d173);
	nor (d266, d99, d164);
	xor (d267, d139, d153);
	and (d268, d114, d159);
	not (d269, d63);
	assign f1 = d223;
	assign f2 = d238;
	assign f3 = d255;
	assign f4 = d226;
	assign f5 = d205;
	assign f6 = d190;
	assign f7 = d195;
	assign f8 = d218;
	assign f9 = d201;
	assign f10 = d184;
	assign f11 = d187;
	assign f12 = d232;
	assign f13 = d253;
	assign f14 = d213;
	assign f15 = d194;
	assign f16 = d224;
	assign f17 = d222;
	assign f18 = d185;
	assign f19 = d256;
endmodule
