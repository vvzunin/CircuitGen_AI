module CCGRCG64( x0, x1, x2, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15 );

	input x0, x1, x2;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265;

	buf (d1, x2);
	nor (d2, x0, x1);
	xor (d3, x1, x2);
	and (d4, x1);
	or (d5, x0, x1);
	and (d6, x0, x1);
	nor (d7, x1, x2);
	xnor (d8, x0, x2);
	nand (d9, x2);
	buf (d10, x1);
	xnor (d11, x1, x2);
	and (d12, x1, x2);
	nand (d13, x0, x2);
	nor (d14, x0, x2);
	buf (d15, x0);
	nor (d16, x1);
	nor (d17, x0);
	or (d18, x1, x2);
	nand (d19, x0, x1);
	and (d20, x1, x2);
	and (d21, x0, x2);
	xor (d22, x0, x2);
	xor (d23, x0, x1);
	or (d24, x2);
	nand (d25, x1, x2);
	not (d26, x1);
	xnor (d27, x0, x1);
	not (d28, x2);
	or (d29, x0);
	and (d30, x0, x1);
	and (d31, x2);
	and (d32, x0, x2);
	and (d33, x0);
	or (d34, x1);
	xnor (d35, x0);
	nand (d36, x0, x2);
	nor (d37, x0, x2);
	not (d38, x0);
	xnor (d39, x0, x2);
	xor (d40, x2);
	xor (d41, x0);
	or (d42, x0, x2);
	xor (d43, x0, x1);
	xor (d44, d2, d6);
	and (d45, d37, d42);
	xnor (d46, d1, d40);
	buf (d47, d26);
	or (d48, d3, d5);
	not (d49, d20);
	xor (d50, d26, d35);
	xnor (d51, d36, d39);
	buf (d52, d24);
	buf (d53, d43);
	nand (d54, d29, d35);
	nand (d55, d8, d34);
	and (d56, d19, d23);
	buf (d57, d5);
	xnor (d58, d17, d28);
	or (d59, d10, d15);
	nor (d60, d1, d40);
	not (d61, d3);
	xnor (d62, d5, d7);
	buf (d63, d27);
	and (d64, d9, d23);
	xnor (d65, d5);
	not (d66, d25);
	xor (d67, d3, d10);
	buf (d68, d8);
	or (d69, d20, d33);
	or (d70, d13, d16);
	nor (d71, d8, d33);
	not (d72, d19);
	nand (d73, d4, d42);
	buf (d74, d32);
	xnor (d75, d36, d41);
	nand (d76, d18, d29);
	xor (d77, d35, d36);
	xnor (d78, d10, d34);
	or (d79, d1, d14);
	and (d80, d3, d34);
	xnor (d81, d24, d26);
	and (d82, d7, d39);
	xor (d83, d10, d32);
	not (d84, d2);
	xnor (d85, d51, d63);
	buf (d86, d6);
	nand (d87, d49, d53);
	and (d88, d64, d70);
	xor (d89, d50, d60);
	xnor (d90, d44, d82);
	nor (d91, d65, d68);
	nor (d92, d68, d74);
	buf (d93, d4);
	nand (d94, d74, d81);
	buf (d95, d25);
	nand (d96, d49, d70);
	xor (d97, d46, d55);
	xor (d98, d60, d75);
	not (d99, d15);
	or (d100, d44, d56);
	nand (d101, d50, d69);
	or (d102, d45, d71);
	xnor (d103, d56, d59);
	or (d104, d58, d70);
	or (d105, d69, d76);
	or (d106, d51, d74);
	and (d107, d65, d75);
	and (d108, d68, d83);
	nor (d109, d44, d56);
	nor (d110, d61, d66);
	buf (d111, d1);
	nor (d112, d50, d59);
	xor (d113, d57, d82);
	not (d114, d30);
	or (d115, d71, d75);
	or (d116, d56, d70);
	and (d117, d67, d80);
	xor (d118, d71, d73);
	nor (d119, d60, d69);
	not (d120, d76);
	not (d121, d55);
	and (d122, d52, d81);
	nor (d123, d51, d71);
	or (d124, d58, d68);
	or (d125, d48, d49);
	xnor (d126, d61, d73);
	xor (d127, d44, d70);
	nor (d128, d71, d74);
	or (d129, d51, d75);
	and (d130, d73, d80);
	xnor (d131, d48, d55);
	nand (d132, d53, d57);
	not (d133, d47);
	and (d134, d79, d81);
	xor (d135, d45, d66);
	or (d136, d50, d59);
	xnor (d137, d63, d76);
	xnor (d138, d61, d66);
	xor (d139, d58, d80);
	nor (d140, d65, d69);
	or (d141, d47, d62);
	xor (d142, d45, d83);
	or (d143, d44, d66);
	buf (d144, d23);
	and (d145, d56, d59);
	xnor (d146, d52, d60);
	xor (d147, d45, d73);
	xor (d148, d52, d79);
	not (d149, d21);
	and (d150, d44, d67);
	not (d151, d18);
	xor (d152, d49, d58);
	not (d153, d41);
	nor (d154, d71, d82);
	buf (d155, d63);
	nand (d156, d45, d47);
	or (d157, d74, d84);
	nor (d158, d58, d65);
	xnor (d159, d65, d79);
	and (d160, d45, d47);
	nand (d161, d57, d72);
	xnor (d162, d47, d57);
	nor (d163, d54, d80);
	or (d164, d62, d84);
	nor (d165, d68, d69);
	nand (d166, d60, d82);
	not (d167, d56);
	and (d168, d51, d74);
	nand (d169, d48, d53);
	buf (d170, d48);
	nor (d171, d55, d73);
	nand (d172, d61, d81);
	nand (d173, d65, d67);
	buf (d174, d19);
	or (d175, d55, d58);
	xor (d176, d53, d75);
	xor (d177, d58, d82);
	xnor (d178, d55, d80);
	xnor (d179, d70, d71);
	xor (d180, d53, d59);
	nand (d181, d160, d177);
	xor (d182, d114, d132);
	nor (d183, d122, d134);
	or (d184, d98, d115);
	xor (d185, d98, d148);
	xor (d186, d105, d139);
	or (d187, d132, d153);
	xor (d188, d119, d134);
	nor (d189, d171, d179);
	xnor (d190, d152, d153);
	nand (d191, d86, d116);
	xor (d192, d115, d145);
	nand (d193, d105, d122);
	not (d194, d164);
	nand (d195, d123, d151);
	or (d196, d96, d123);
	nor (d197, d171, d178);
	xor (d198, d125, d135);
	nand (d199, d87, d120);
	nor (d200, d110, d169);
	or (d201, d105, d149);
	or (d202, d114, d141);
	and (d203, d143, d164);
	or (d204, d112, d172);
	xor (d205, d85, d174);
	xnor (d206, d86, d133);
	nor (d207, d89, d161);
	not (d208, d79);
	or (d209, d94, d179);
	and (d210, d94, d106);
	nand (d211, d119, d130);
	and (d212, d163, d169);
	nand (d213, d86, d128);
	xnor (d214, d105, d124);
	not (d215, d171);
	nand (d216, d86, d168);
	nand (d217, d128, d152);
	nor (d218, d138, d159);
	not (d219, d113);
	nand (d220, d121, d124);
	xor (d221, d137, d164);
	xnor (d222, d99, d167);
	xor (d223, d169, d172);
	buf (d224, d167);
	buf (d225, d103);
	xor (d226, d104, d148);
	xnor (d227, d119, d142);
	or (d228, d116, d169);
	xor (d229, d107, d119);
	or (d230, d98, d167);
	not (d231, d102);
	not (d232, d152);
	and (d233, d114, d155);
	xor (d234, d173, d178);
	xor (d235, d85, d174);
	nand (d236, d95, d120);
	nor (d237, d133, d139);
	nor (d238, d170, d178);
	nor (d239, d102, d167);
	nand (d240, d88, d99);
	xnor (d241, d95, d164);
	buf (d242, d118);
	xor (d243, d140, d161);
	and (d244, d99, d177);
	or (d245, d123, d161);
	and (d246, d130, d178);
	or (d247, d160, d171);
	and (d248, d86, d141);
	xor (d249, d91, d177);
	xnor (d250, d140, d165);
	xor (d251, d86, d157);
	nor (d252, d116, d176);
	and (d253, d100, d144);
	xor (d254, d135, d152);
	not (d255, d125);
	not (d256, d163);
	and (d257, d171, d177);
	not (d258, d34);
	and (d259, d154, d180);
	xor (d260, d123, d164);
	buf (d261, d64);
	xnor (d262, d95, d98);
	not (d263, d103);
	or (d264, d111, d118);
	nor (d265, d88, d146);
	assign f1 = d207;
	assign f2 = d182;
	assign f3 = d240;
	assign f4 = d200;
	assign f5 = d251;
	assign f6 = d229;
	assign f7 = d260;
	assign f8 = d212;
	assign f9 = d214;
	assign f10 = d264;
	assign f11 = d229;
	assign f12 = d237;
	assign f13 = d229;
	assign f14 = d234;
	assign f15 = d185;
endmodule
