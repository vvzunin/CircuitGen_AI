module CCGRCG94( x0, x1, x2, x3, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11 );

	input x0, x1, x2, x3;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264;

	or (d1, x0, x2);
	xnor (d2, x0, x2);
	and (d3, x2);
	xnor (d4, x1);
	nand (d5, x0, x3);
	buf (d6, x3);
	and (d7, x0, x2);
	and (d8, x1, x2);
	not (d9, x0);
	nand (d10, x1, x3);
	and (d11, x0, x3);
	and (d12, x3);
	xnor (d13, x0, x3);
	buf (d14, x0);
	not (d15, x2);
	or (d16, x0, x3);
	xor (d17, x0, x1);
	and (d18, x1, x2);
	nand (d19, x0, x1);
	not (d20, d13);
	nor (d21, d9, d14);
	nor (d22, d11, d18);
	nor (d23, d2, d16);
	not (d24, d10);
	buf (d25, d4);
	xnor (d26, d1, d4);
	buf (d27, d1);
	nor (d28, d7, d15);
	xnor (d29, d9, d17);
	xor (d30, d1, d4);
	buf (d31, d13);
	or (d32, d5, d10);
	or (d33, d13, d14);
	or (d34, d6, d14);
	xnor (d35, d18);
	xnor (d36, d2, d17);
	not (d37, d12);
	and (d38, d13, d17);
	buf (d39, d5);
	and (d40, d8, d16);
	nand (d41, d12, d18);
	and (d42, d7, d12);
	xnor (d43, d12, d17);
	xnor (d44, d11, d15);
	nor (d45, d4, d5);
	xnor (d46, d8, d14);
	nand (d47, d1, d12);
	not (d48, d5);
	and (d49, d16, d18);
	not (d50, x3);
	xor (d51, d8, d16);
	buf (d52, d16);
	nor (d53, d4, d11);
	not (d54, d9);
	nor (d55, d12, d18);
	xor (d56, d1, d15);
	nor (d57, d6, d9);
	and (d58, d14, d16);
	not (d59, d3);
	nor (d60, d8, d19);
	xor (d61, d2, d15);
	nor (d62, d10, d14);
	nand (d63, d12, d19);
	xor (d64, d1, d19);
	xor (d65, d9, d18);
	xnor (d66, d5, d11);
	xor (d67, d1, d7);
	or (d68, d7, d9);
	nand (d69, d2, d12);
	buf (d70, d9);
	xor (d71, d4, d19);
	nor (d72, d13, d17);
	buf (d73, d11);
	xor (d74, d10, d13);
	or (d75, d8, d11);
	nand (d76, d3, d17);
	and (d77, d1, d19);
	xnor (d78, d3, d11);
	xnor (d79, d4, d19);
	not (d80, d6);
	and (d81, d6, d9);
	or (d82, d7, d15);
	and (d83, d8, d18);
	not (d84, d4);
	nor (d85, d7, d9);
	nor (d86, d16);
	xnor (d87, d9);
	xor (d88, d4, d6);
	and (d89, d1);
	nor (d90, d18);
	nand (d91, d1, d15);
	or (d92, d2, d15);
	and (d93, d17, d19);
	xor (d94, d3);
	and (d95, d8, d17);
	xnor (d96, d1);
	or (d97, d7);
	nand (d98, d1, d13);
	nand (d99, d53, d87);
	nor (d100, d24, d50);
	xnor (d101, d78, d90);
	xnor (d102, d49, d81);
	or (d103, d24, d25);
	nand (d104, d46, d58);
	nor (d105, d41, d61);
	not (d106, d80);
	nand (d107, d87, d98);
	not (d108, d69);
	nand (d109, d50, d93);
	or (d110, d41, d61);
	not (d111, d35);
	xnor (d112, d21, d91);
	nand (d113, d60, d73);
	xnor (d114, d50, d93);
	not (d115, d50);
	buf (d116, d92);
	or (d117, d22, d80);
	nand (d118, d85, d89);
	buf (d119, d95);
	or (d120, d66, d93);
	xnor (d121, d22, d89);
	nor (d122, d27, d69);
	nor (d123, d61, d93);
	buf (d124, x2);
	buf (d125, d2);
	buf (d126, d76);
	nand (d127, d51, d53);
	nand (d128, d72, d86);
	buf (d129, d35);
	xnor (d130, d23, d66);
	nand (d131, d75, d89);
	xnor (d132, d20, d44);
	not (d133, d55);
	or (d134, d24, d39);
	nand (d135, d33, d96);
	not (d136, d95);
	xnor (d137, d20, d46);
	xor (d138, d74, d84);
	and (d139, d52, d66);
	xnor (d140, d21, d84);
	xnor (d141, d62, d73);
	not (d142, d28);
	not (d143, d73);
	nor (d144, d26, d97);
	nor (d145, d25, d53);
	and (d146, d60, d69);
	xnor (d147, d38, d53);
	xnor (d148, d25, d34);
	not (d149, d76);
	or (d150, d34, d43);
	or (d151, d44, d82);
	buf (d152, d53);
	and (d153, d30, d79);
	nor (d154, d92, d98);
	and (d155, d30, d68);
	and (d156, d49, d69);
	xnor (d157, d21, d83);
	nand (d158, d42, d46);
	nor (d159, d30, d50);
	xor (d160, d66, d79);
	xnor (d161, d20, d55);
	xnor (d162, d28, d97);
	not (d163, d67);
	and (d164, d26, d74);
	nand (d165, d20, d70);
	or (d166, d33, d85);
	and (d167, d58, d88);
	buf (d168, d25);
	xor (d169, d48, d58);
	and (d170, d47, d68);
	nand (d171, d55, d71);
	xor (d172, d50, d51);
	nor (d173, d63, d77);
	xor (d174, d20, d36);
	or (d175, d26, d66);
	and (d176, d40, d52);
	nor (d177, d31, d36);
	buf (d178, d28);
	buf (d179, d72);
	and (d180, d23, d66);
	nor (d181, d81, d83);
	xnor (d182, d56, d61);
	xnor (d183, d62, d79);
	buf (d184, d51);
	buf (d185, d82);
	xnor (d186, d86, d87);
	not (d187, d154);
	xnor (d188, d144, d169);
	or (d189, d168, d182);
	nand (d190, d100, d112);
	nor (d191, d111, d166);
	not (d192, d46);
	not (d193, d155);
	xnor (d194, d112, d177);
	xnor (d195, d122, d148);
	nor (d196, d130, d183);
	nor (d197, d129, d172);
	not (d198, d104);
	nor (d199, d197, d198);
	xnor (d200, d188, d195);
	xor (d201, d187, d194);
	nor (d202, d198);
	xor (d203, d194, d197);
	not (d204, d54);
	buf (d205, d195);
	not (d206, d161);
	or (d207, d189, d195);
	and (d208, d194, d197);
	nor (d209, d189, d194);
	and (d210, d188, d192);
	buf (d211, d131);
	or (d212, d191, d192);
	nor (d213, d191, d195);
	nand (d214, d189, d191);
	nand (d215, d196);
	xnor (d216, d191, d196);
	or (d217, d193, d198);
	buf (d218, d166);
	nor (d219, d189, d194);
	xnor (d220, d187, d189);
	or (d221, d192, d197);
	nor (d222, d188, d195);
	buf (d223, d81);
	xnor (d224, d191, d194);
	or (d225, d189, d198);
	and (d226, d188, d191);
	xor (d227, d196, d198);
	not (d228, d65);
	not (d229, d100);
	or (d230, d189, d191);
	and (d231, d189, d198);
	not (d232, d153);
	or (d233, d191, d194);
	buf (d234, d38);
	and (d235, d195, d196);
	xnor (d236, d187, d196);
	xor (d237, d187, d189);
	and (d238, d192, d193);
	xor (d239, d192, d194);
	xor (d240, d196, d198);
	xor (d241, d188, d189);
	buf (d242, d193);
	and (d243, d188, d190);
	buf (d244, d36);
	buf (d245, d175);
	or (d246, d195, d197);
	nand (d247, d191, d198);
	xor (d248, d192, d194);
	nand (d249, d189, d196);
	or (d250, d188, d196);
	nand (d251, d195, d197);
	nand (d252, d190, d191);
	not (d253, d170);
	or (d254, d187, d197);
	or (d255, d188, d189);
	xor (d256, d192, d198);
	not (d257, d145);
	xnor (d258, d193, d196);
	and (d259, d189, d192);
	nand (d260, d192, d196);
	nor (d261, d187, d195);
	nand (d262, d189, d193);
	xnor (d263, d191, d197);
	and (d264, d193, d198);
	assign f1 = d245;
	assign f2 = d264;
	assign f3 = d201;
	assign f4 = d238;
	assign f5 = d211;
	assign f6 = d210;
	assign f7 = d255;
	assign f8 = d244;
	assign f9 = d210;
	assign f10 = d260;
	assign f11 = d209;
endmodule
