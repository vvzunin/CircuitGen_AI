module CCGRCG179( x0, x1, x2, x3, x4, x5, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15 );

	input x0, x1, x2, x3, x4, x5;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169;

	not (d1, x4);
	buf (d2, x2);
	xor (d3, x0);
	or (d4, x2, x3);
	nand (d5, x0, x5);
	or (d6, x1, x5);
	not (d7, x3);
	xor (d8, x0, x3);
	or (d9, x1, x5);
	xor (d10, x3, x4);
	nor (d11, x0, x3);
	xor (d12, x4);
	nand (d13, x0, x4);
	and (d14, x5);
	not (d15, x1);
	xnor (d16, x3, x5);
	buf (d17, x3);
	or (d18, x4);
	xor (d19, x0, x3);
	nor (d20, x1, x3);
	xnor (d21, x1);
	nand (d22, x3, x4);
	nor (d23, x1);
	xnor (d24, x0, x2);
	and (d25, x0, x1);
	nand (d26, x3, x4);
	nor (d27, x3, x4);
	xor (d28, x4, x5);
	and (d29, x2, x5);
	xor (d30, x2, x3);
	xor (d31, x2, x5);
	not (d32, x2);
	buf (d33, x0);
	xnor (d34, x0, x4);
	xnor (d35, x1, x2);
	buf (d36, x1);
	and (d37, x3, x4);
	nand (d38, x3, x5);
	buf (d39, x5);
	nand (d40, x0, x2);
	xor (d41, x2, x4);
	nand (d42, x2, x3);
	xnor (d43, x0, x4);
	and (d44, x1, x5);
	or (d45, x2);
	nor (d46, x0, x1);
	or (d47, x0, x1);
	nor (d48, x3, x4);
	xnor (d49, x0, x2);
	nand (d50, x1, x2);
	xnor (d51, x0, x3);
	or (d52, x0, x4);
	and (d53, x1, x4);
	nand (d54, x0, x2);
	or (d55, x1, x3);
	nand (d56, x1);
	nand (d57, x1, x5);
	and (d58, x4, x5);
	buf (d59, x4);
	nor (d60, x2, x5);
	nand (d61, x3, x5);
	nor (d62, x1, x5);
	or (d63, x1, x2);
	nand (d64, x2);
	xor (d65, d9, d48);
	and (d66, d51, d64);
	not (d67, d61);
	or (d68, d11, d43);
	or (d69, d18, d27);
	nor (d70, d22, d49);
	not (d71, d38);
	nor (d72, d27, d34);
	xnor (d73, d20, d53);
	buf (d74, d37);
	nor (d75, d3, d13);
	or (d76, d29, d47);
	nand (d77, d7, d36);
	nor (d78, d12, d42);
	buf (d79, d48);
	nand (d80, d13, d63);
	or (d81, d69, d73);
	or (d82, d66, d77);
	xor (d83, d65, d80);
	nand (d84, d71, d76);
	buf (d85, d26);
	buf (d86, d41);
	buf (d87, d47);
	buf (d88, d4);
	nand (d89, d74, d77);
	not (d90, d14);
	not (d91, d59);
	buf (d92, d45);
	nor (d93, d73, d80);
	or (d94, d68, d79);
	xor (d95, d69, d79);
	and (d96, d68, d75);
	nor (d97, d72, d79);
	nand (d98, d68, d77);
	nand (d99, d78, d80);
	buf (d100, d64);
	and (d101, d69, d75);
	or (d102, d76, d78);
	or (d103, d70, d76);
	or (d104, d65, d73);
	nor (d105, d70, d71);
	and (d106, d76);
	xnor (d107, d65, d71);
	xnor (d108, d79, d80);
	not (d109, d54);
	xor (d110, d80);
	or (d111, d69, d77);
	or (d112, d73, d76);
	xnor (d113, d72, d78);
	xor (d114, d76, d80);
	not (d115, d33);
	nand (d116, d65, d73);
	buf (d117, d53);
	or (d118, d72, d74);
	or (d119, d73, d77);
	not (d120, d56);
	nor (d121, d75, d79);
	buf (d122, d35);
	nor (d123, d74, d77);
	xnor (d124, d67, d71);
	nor (d125, d75, d77);
	or (d126, d72, d73);
	nand (d127, d68, d69);
	not (d128, d4);
	and (d129, d70, d74);
	or (d130, d78);
	xor (d131, d71, d73);
	xnor (d132, d73, d76);
	not (d133, d43);
	buf (d134, d44);
	nand (d135, d73, d74);
	xor (d136, d67, d78);
	xor (d137, d68, d79);
	and (d138, d75, d78);
	not (d139, d44);
	nor (d140, d67, d77);
	nor (d141, d65, d80);
	buf (d142, d78);
	and (d143, d73);
	xnor (d144, d71, d75);
	and (d145, d68, d78);
	not (d146, d46);
	xor (d147, d79, d80);
	xor (d148, d66, d67);
	nor (d149, d78, d80);
	xor (d150, d66, d69);
	or (d151, d68, d73);
	nor (d152, d69, d76);
	xor (d153, d69, d80);
	not (d154, d12);
	or (d155, d77, d79);
	not (d156, d7);
	nor (d157, d65, d77);
	xnor (d158, d77, d79);
	not (d159, d50);
	not (d160, d75);
	or (d161, d71, d76);
	nor (d162, d66, d79);
	buf (d163, d7);
	nor (d164, d70, d72);
	nand (d165, d76, d79);
	xnor (d166, d73, d80);
	not (d167, d15);
	and (d168, d72, d76);
	buf (d169, d63);
	assign f1 = d134;
	assign f2 = d135;
	assign f3 = d110;
	assign f4 = d104;
	assign f5 = d144;
	assign f6 = d164;
	assign f7 = d90;
	assign f8 = d94;
	assign f9 = d149;
	assign f10 = d104;
	assign f11 = d134;
	assign f12 = d148;
	assign f13 = d161;
	assign f14 = d158;
	assign f15 = d153;
endmodule
