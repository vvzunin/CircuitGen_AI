module CCGRCG98( x0, x1, x2, x3, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13 );

	input x0, x1, x2, x3;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314, d315, d316, d317, d318, d319, d320, d321, d322, d323, d324, d325, d326, d327, d328, d329, d330, d331, d332, d333, d334, d335, d336, d337, d338, d339, d340, d341, d342, d343, d344, d345, d346, d347, d348, d349, d350, d351, d352, d353, d354, d355, d356, d357, d358, d359, d360, d361, d362, d363, d364, d365, d366, d367, d368, d369, d370, d371, d372, d373, d374, d375, d376, d377, d378, d379, d380, d381, d382, d383, d384, d385, d386, d387, d388, d389, d390, d391, d392, d393, d394, d395, d396, d397, d398, d399, d400, d401, d402, d403, d404, d405, d406, d407, d408, d409, d410, d411, d412, d413, d414, d415, d416, d417, d418, d419, d420, d421, d422, d423, d424, d425, d426, d427, d428, d429, d430, d431, d432, d433, d434, d435, d436, d437, d438, d439, d440, d441, d442, d443, d444, d445, d446, d447, d448, d449, d450, d451, d452, d453, d454;

	xnor (d1, x0, x2);
	not (d2, x3);
	buf (d3, x1);
	xor (d4, x1, x3);
	buf (d5, x3);
	not (d6, x2);
	buf (d7, x2);
	xnor (d8, x0, x1);
	nand (d9, x2, x3);
	xor (d10, x0, x3);
	nor (d11, x2);
	or (d12, x2, x3);
	nor (d13, x1);
	buf (d14, x0);
	and (d15, x2, x3);
	and (d16, x0, x3);
	or (d17, x1, x3);
	or (d18, x0, x2);
	nand (d19, x1, x2);
	xnor (d20, x1, x3);
	xnor (d21, x2);
	xor (d22, x0, x2);
	or (d23, x0);
	xnor (d24, x2, x3);
	xor (d25, x0, x1);
	xnor (d26, x1, x2);
	xor (d27, d6, d7);
	not (d28, d23);
	xnor (d29, d15, d26);
	nor (d30, d20);
	not (d31, x1);
	buf (d32, d13);
	and (d33, d11, d20);
	xor (d34, d13, d26);
	or (d35, d5, d11);
	buf (d36, d14);
	buf (d37, d23);
	nand (d38, d9, d22);
	or (d39, d12, d13);
	nand (d40, d2, d17);
	nand (d41, d18, d19);
	nand (d42, d7, d12);
	xor (d43, d20, d25);
	and (d44, d3, d17);
	and (d45, d7, d23);
	xnor (d46, d16, d20);
	nor (d47, d3, d22);
	xor (d48, d3);
	xnor (d49, d5, d17);
	nor (d50, d6, d23);
	not (d51, d18);
	nor (d52, d1, d19);
	nand (d53, d4, d26);
	xnor (d54, d7, d8);
	xor (d55, d1, d26);
	and (d56, d12, d24);
	and (d57, d4, d6);
	and (d58, d1, d21);
	nor (d59, d5, d16);
	nor (d60, d14, d24);
	not (d61, d20);
	nand (d62, d18, d20);
	not (d63, d11);
	not (d64, d19);
	xnor (d65, d8, d12);
	nand (d66, d12, d21);
	nor (d67, d7, d18);
	nor (d68, d9, d18);
	or (d69, d22, d26);
	nor (d70, d13, d15);
	nor (d71, d8, d25);
	not (d72, d16);
	nand (d73, d11, d15);
	xor (d74, d6, d23);
	xnor (d75, d3, d23);
	xnor (d76, d1, d15);
	nand (d77, d8, d14);
	xor (d78, d7, d18);
	xor (d79, d11, d20);
	nand (d80, d19, d24);
	and (d81, d9, d10);
	nor (d82, d11, d15);
	nand (d83, d2, d14);
	and (d84, d3, d14);
	xnor (d85, d4, d10);
	nor (d86, d13, d16);
	not (d87, d1);
	or (d88, d3, d19);
	and (d89, d14, d21);
	not (d90, d13);
	xnor (d91, d1, d2);
	xnor (d92, d11, d12);
	xor (d93, d10, d22);
	xnor (d94, d3);
	not (d95, d26);
	and (d96, d17, d26);
	nor (d97, d18, d20);
	or (d98, d19, d25);
	xor (d99, d2, d7);
	and (d100, d5, d13);
	nor (d101, d32, d87);
	xnor (d102, d56, d91);
	nand (d103, d40, d82);
	xnor (d104, d55, d90);
	xnor (d105, d45, d89);
	buf (d106, d15);
	nand (d107, d32, d91);
	buf (d108, d92);
	or (d109, d42, d52);
	not (d110, d45);
	nor (d111, d74, d96);
	or (d112, d48, d69);
	nand (d113, d36, d59);
	buf (d114, d17);
	and (d115, d79, d83);
	buf (d116, d38);
	not (d117, d12);
	nand (d118, d53, d73);
	buf (d119, d96);
	and (d120, d85, d87);
	xnor (d121, d65, d88);
	and (d122, d91, d92);
	xnor (d123, d54, d94);
	xor (d124, d28, d94);
	xnor (d125, d37, d76);
	and (d126, d77, d84);
	xnor (d127, d64, d79);
	nand (d128, d78, d98);
	xor (d129, d80, d100);
	not (d130, d87);
	nor (d131, d72, d79);
	xor (d132, d70, d94);
	nand (d133, d72, d84);
	buf (d134, d46);
	and (d135, d35, d49);
	or (d136, d48, d88);
	xor (d137, d92, d100);
	not (d138, d6);
	buf (d139, d9);
	nor (d140, d73, d90);
	and (d141, d33, d67);
	buf (d142, d40);
	or (d143, d31, d40);
	buf (d144, d54);
	nor (d145, d44, d47);
	buf (d146, d97);
	not (d147, d15);
	or (d148, d68, d94);
	buf (d149, d52);
	buf (d150, d30);
	xor (d151, d66, d71);
	and (d152, d53, d69);
	or (d153, d46, d79);
	and (d154, d40, d98);
	buf (d155, d10);
	nand (d156, d76, d80);
	or (d157, d44, d78);
	and (d158, d28, d40);
	nand (d159, d45, d96);
	nor (d160, d63, d97);
	and (d161, d53, d73);
	nand (d162, d145, d148);
	or (d163, d104, d127);
	buf (d164, d50);
	buf (d165, d36);
	buf (d166, d31);
	buf (d167, d139);
	not (d168, d107);
	buf (d169, d18);
	and (d170, d125, d140);
	or (d171, d138);
	nand (d172, d108, d145);
	xor (d173, d135, d144);
	and (d174, d117, d155);
	nand (d175, d134, d158);
	nor (d176, d113, d139);
	not (d177, d62);
	xnor (d178, d102, d115);
	buf (d179, d94);
	nor (d180, d122, d139);
	xor (d181, d125, d138);
	nand (d182, d151, d158);
	nand (d183, d108, d110);
	nand (d184, d140, d150);
	or (d185, d114, d157);
	and (d186, d115, d123);
	and (d187, d116, d140);
	xnor (d188, d108, d134);
	buf (d189, d76);
	nand (d190, d102, d151);
	and (d191, d149, d154);
	nor (d192, d119, d150);
	or (d193, d106, d115);
	nor (d194, d115, d158);
	and (d195, d112, d134);
	xnor (d196, d105, d145);
	xor (d197, d122, d153);
	or (d198, d104, d122);
	not (d199, d75);
	xnor (d200, d116, d159);
	or (d201, d119, d157);
	and (d202, d140, d158);
	xor (d203, d135, d157);
	or (d204, d150, d151);
	nand (d205, d146, d152);
	not (d206, d117);
	buf (d207, d69);
	xor (d208, d194, d195);
	nand (d209, d176, d199);
	or (d210, d173, d185);
	and (d211, d192, d196);
	xor (d212, d176, d203);
	not (d213, d30);
	xor (d214, d198, d199);
	nand (d215, d178, d200);
	and (d216, d175, d205);
	nand (d217, d171, d197);
	xnor (d218, d178, d184);
	not (d219, d82);
	xor (d220, d176, d203);
	nand (d221, d169, d182);
	or (d222, d165, d203);
	nor (d223, d163, d205);
	not (d224, d132);
	nor (d225, d194);
	not (d226, d71);
	or (d227, d162, d165);
	xnor (d228, d184, d190);
	nand (d229, d195, d200);
	xor (d230, d175, d195);
	xor (d231, d184, d190);
	buf (d232, d107);
	buf (d233, d157);
	or (d234, d176, d188);
	nor (d235, d174, d198);
	or (d236, d187);
	buf (d237, d111);
	or (d238, d172, d206);
	and (d239, d163, d181);
	or (d240, d186, d199);
	nand (d241, d170, d197);
	nand (d242, d175, d188);
	or (d243, d164, d183);
	buf (d244, d187);
	buf (d245, d180);
	and (d246, d176, d184);
	or (d247, d171, d197);
	nor (d248, d178, d205);
	and (d249, d171, d207);
	nand (d250, d162, d169);
	buf (d251, d80);
	buf (d252, d86);
	xor (d253, d191, d193);
	not (d254, d105);
	xor (d255, d173, d176);
	nand (d256, d166, d173);
	nand (d257, d163, d180);
	or (d258, d173, d191);
	xor (d259, d189, d207);
	nor (d260, d162, d192);
	xnor (d261, d166, d186);
	nor (d262, d186, d195);
	buf (d263, d88);
	xor (d264, d173, d192);
	buf (d265, d148);
	xor (d266, d196, d197);
	and (d267, d191, d194);
	and (d268, d184, d195);
	nor (d269, d171, d201);
	nor (d270, d163, d198);
	or (d271, d187, d206);
	nand (d272, d189);
	xor (d273, d165, d196);
	not (d274, d60);
	and (d275, d168, d189);
	xor (d276, d184, d205);
	buf (d277, d199);
	and (d278, d166, d195);
	xnor (d279, d184, d199);
	xor (d280, d166, d192);
	nand (d281, d169, d172);
	xor (d282, d177, d179);
	nand (d283, d170, d204);
	xnor (d284, d167, d204);
	buf (d285, d43);
	not (d286, d92);
	xor (d287, d179, d205);
	xnor (d288, d194, d195);
	or (d289, d190, d202);
	not (d290, d43);
	not (d291, d180);
	xnor (d292, d175, d201);
	nor (d293, d210, d244);
	xnor (d294, d236, d291);
	not (d295, d216);
	nand (d296, d219, d281);
	not (d297, d153);
	and (d298, d218, d244);
	not (d299, d198);
	xnor (d300, d249, d281);
	buf (d301, d283);
	not (d302, d122);
	buf (d303, d271);
	buf (d304, d217);
	xor (d305, d254, d292);
	nor (d306, d223, d251);
	buf (d307, d2);
	or (d308, d221, d251);
	xor (d309, d228, d289);
	not (d310, d176);
	and (d311, d237, d240);
	nor (d312, d273, d277);
	xor (d313, d229, d239);
	xor (d314, d283, d288);
	not (d315, d191);
	or (d316, d263, d291);
	and (d317, d224, d238);
	xnor (d318, d282, d287);
	xor (d319, d210, d266);
	and (d320, d294, d314);
	buf (d321, d12);
	not (d322, d115);
	nor (d323, d305, d317);
	xnor (d324, d305, d316);
	xnor (d325, d293, d296);
	nor (d326, d302, d305);
	xor (d327, d297, d307);
	nor (d328, d296, d304);
	and (d329, d300, d317);
	xnor (d330, d303, d308);
	or (d331, d294, d310);
	xor (d332, d300, d306);
	xor (d333, d303, d310);
	nor (d334, d296, d298);
	or (d335, d306, d315);
	buf (d336, d6);
	nand (d337, d299, d305);
	not (d338, d183);
	not (d339, d101);
	buf (d340, d45);
	nand (d341, d313, d314);
	or (d342, d300, d305);
	or (d343, d313, d319);
	or (d344, d306, d312);
	nand (d345, d303, d317);
	not (d346, d61);
	nand (d347, d293, d316);
	and (d348, d305, d306);
	xnor (d349, d294, d313);
	xor (d350, d293, d294);
	nor (d351, d301, d307);
	or (d352, d309, d315);
	xnor (d353, d305, d312);
	or (d354, d309, d311);
	nor (d355, d306, d316);
	nor (d356, d294, d299);
	nand (d357, d304, d317);
	nand (d358, d313, d319);
	and (d359, d304, d314);
	nand (d360, d293, d301);
	nand (d361, d313, d317);
	and (d362, d296, d309);
	and (d363, d307, d316);
	xor (d364, d297, d304);
	nor (d365, d296, d308);
	buf (d366, d42);
	and (d367, d295, d298);
	and (d368, d311, d319);
	or (d369, d300, d309);
	nor (d370, d306, d313);
	xnor (d371, d301, d303);
	or (d372, d303, d307);
	buf (d373, d252);
	buf (d374, d213);
	nand (d375, d358, d367);
	not (d376, d47);
	buf (d377, d363);
	xnor (d378, d336, d369);
	not (d379, d257);
	xnor (d380, d350, d364);
	xor (d381, d321, d346);
	or (d382, d337, d368);
	nand (d383, d342, d355);
	buf (d384, d165);
	nand (d385, d341, d368);
	or (d386, d345, d349);
	or (d387, d345);
	and (d388, d354, d361);
	xor (d389, d336, d362);
	xnor (d390, d332, d356);
	nand (d391, d353, d367);
	nor (d392, d338, d340);
	or (d393, d338, d370);
	xor (d394, d331, d358);
	nor (d395, d323, d337);
	xor (d396, d358, d371);
	xnor (d397, d355, d372);
	nand (d398, d344, d357);
	buf (d399, d248);
	xnor (d400, d337, d349);
	xnor (d401, d321, d351);
	not (d402, d239);
	and (d403, d321, d359);
	or (d404, d320, d340);
	nand (d405, d331, d366);
	nand (d406, d320, d358);
	xor (d407, d326);
	xnor (d408, d329, d357);
	xor (d409, d335, d347);
	nor (d410, d341, d358);
	not (d411, d221);
	buf (d412, d70);
	xor (d413, d383, d385);
	buf (d414, d336);
	nand (d415, d377, d386);
	and (d416, d388, d399);
	nand (d417, d393, d395);
	nand (d418, d380, d383);
	nor (d419, d381, d399);
	and (d420, d397);
	or (d421, d383, d400);
	buf (d422, d172);
	or (d423, d378, d381);
	nand (d424, d388, d391);
	xor (d425, d406, d410);
	buf (d426, d196);
	xor (d427, d381, d396);
	or (d428, d373, d409);
	nor (d429, d393, d407);
	or (d430, d392, d399);
	xor (d431, d375, d380);
	nor (d432, d388, d393);
	and (d433, d378, d404);
	nor (d434, d388, d407);
	xor (d435, d390, d396);
	nor (d436, d395, d402);
	and (d437, d383, d409);
	nand (d438, d373, d379);
	xor (d439, d390, d398);
	nor (d440, d380, d390);
	xor (d441, d398, d409);
	or (d442, d391, d392);
	or (d443, d395, d406);
	nand (d444, d376, d400);
	and (d445, d379, d390);
	xnor (d446, d389, d397);
	nand (d447, d389, d395);
	not (d448, d321);
	not (d449, d83);
	xor (d450, d373, d407);
	or (d451, d387, d407);
	xnor (d452, d388, d399);
	nand (d453, d383, d391);
	nand (d454, d396, d409);
	assign f1 = d414;
	assign f2 = d449;
	assign f3 = d424;
	assign f4 = d415;
	assign f5 = d439;
	assign f6 = d420;
	assign f7 = d440;
	assign f8 = d412;
	assign f9 = d430;
	assign f10 = d431;
	assign f11 = d412;
	assign f12 = d449;
	assign f13 = d427;
endmodule
