module CCGRCG103( x0, x1, x2, x3, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15 );

	input x0, x1, x2, x3;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145;

	and (d1, x0, x1);
	xnor (d2, x0, x2);
	not (d3, x3);
	nor (d4, x0);
	not (d5, x0);
	and (d6, x1, x2);
	and (d7, x2, x3);
	or (d8, x0, x2);
	and (d9, x0, x3);
	not (d10, x2);
	nor (d11, x0, x1);
	nor (d12, x1, x3);
	buf (d13, x2);
	or (d14, x2);
	buf (d15, x0);
	nor (d16, x0, x2);
	xnor (d17, x2, x3);
	or (d18, x0, x1);
	and (d19, x0, x3);
	nor (d20, x1, x2);
	nor (d21, x2);
	nor (d22, x1, x3);
	nand (d23, x0, x1);
	nor (d24, x1);
	nor (d25, x0, x3);
	nor (d26, x3);
	xnor (d27, x0, x1);
	xor (d28, x0, x3);
	buf (d29, x1);
	nor (d30, x2, x3);
	nand (d31, x2, x3);
	xor (d32, x0);
	nor (d33, x2, x3);
	not (d34, x1);
	xor (d35, x1, x3);
	xor (d36, x2, x3);
	or (d37, x0);
	nand (d38, x1, x3);
	nand (d39, x0, x3);
	nor (d40, x0, x2);
	xor (d41, x2, x3);
	buf (d42, x3);
	and (d43, x0);
	nand (d44, x1, x2);
	xnor (d45, x1);
	xor (d46, x1, x3);
	xor (d47, x0, x3);
	xnor (d48, x2, x3);
	and (d49, x3);
	or (d50, x3);
	xor (d51, x1);
	nand (d52, d22, d25);
	xnor (d53, d48);
	xor (d54, d6, d14);
	not (d55, d2);
	not (d56, d13);
	not (d57, d36);
	buf (d58, d26);
	xnor (d59, d15, d35);
	buf (d60, d23);
	xnor (d61, d45, d47);
	not (d62, d35);
	not (d63, d40);
	or (d64, d11, d19);
	and (d65, d41, d42);
	xnor (d66, d26, d33);
	xnor (d67, d10, d46);
	nand (d68, d46, d47);
	nand (d69, d24, d26);
	nand (d70, d1, d24);
	nand (d71, d26, d46);
	xor (d72, d5, d13);
	nand (d73, d7, d13);
	nand (d74, d10, d22);
	xnor (d75, d5, d27);
	xnor (d76, d6, d11);
	xnor (d77, d8, d26);
	xnor (d78, d15, d25);
	and (d79, d16, d35);
	and (d80, d18, d30);
	buf (d81, d47);
	nand (d82, d15, d35);
	nor (d83, d28, d51);
	xor (d84, d35, d50);
	xor (d85, d33, d45);
	nand (d86, d23, d31);
	xnor (d87, d29, d42);
	not (d88, d12);
	xor (d89, d15, d38);
	nor (d90, d1, d32);
	nor (d91, d39, d41);
	xor (d92, d13, d31);
	buf (d93, d49);
	nand (d94, d11, d37);
	or (d95, d24, d32);
	xnor (d96, d6, d18);
	nand (d97, d16, d35);
	xor (d98, d17, d27);
	xnor (d99, d30, d36);
	xor (d100, d3, d42);
	buf (d101, d32);
	xnor (d102, d4, d28);
	nand (d103, d3, d46);
	xnor (d104, d42, d44);
	and (d105, d11, d19);
	xor (d106, d26, d43);
	or (d107, d32, d36);
	and (d108, d26, d29);
	xor (d109, d19, d37);
	xnor (d110, d7, d39);
	or (d111, d11, d51);
	nor (d112, d16, d34);
	xor (d113, d8, d36);
	buf (d114, d22);
	nand (d115, d20, d33);
	or (d116, d42, d51);
	nor (d117, d13, d27);
	or (d118, d2, d29);
	xnor (d119, d34, d37);
	xor (d120, d50);
	not (d121, d37);
	nand (d122, d4, d23);
	nor (d123, d10, d43);
	not (d124, d1);
	xnor (d125, d6, d27);
	xor (d126, d1, d12);
	xnor (d127, d35, d36);
	nand (d128, d11, d20);
	or (d129, d27, d49);
	nor (d130, d21, d23);
	and (d131, d9, d46);
	xor (d132, d36, d47);
	not (d133, d18);
	not (d134, d21);
	nand (d135, d5, d48);
	nor (d136, d20, d26);
	xor (d137, d23, d51);
	and (d138, d20, d36);
	or (d139, d34, d48);
	xnor (d140, d10, d40);
	not (d141, d24);
	xor (d142, d3, d19);
	xor (d143, d19, d47);
	or (d144, d17, d26);
	nor (d145, d48, d51);
	assign f1 = d129;
	assign f2 = d69;
	assign f3 = d79;
	assign f4 = d106;
	assign f5 = d111;
	assign f6 = d85;
	assign f7 = d130;
	assign f8 = d128;
	assign f9 = d128;
	assign f10 = d98;
	assign f11 = d81;
	assign f12 = d126;
	assign f13 = d87;
	assign f14 = d143;
	assign f15 = d62;
endmodule
