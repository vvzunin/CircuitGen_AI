module CCGRCG177( x0, x1, x2, x3, x4, x5, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14 );

	input x0, x1, x2, x3, x4, x5;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314, d315, d316, d317, d318, d319, d320, d321, d322, d323, d324, d325, d326, d327, d328, d329, d330, d331, d332, d333, d334, d335, d336, d337, d338, d339, d340, d341, d342, d343, d344, d345, d346, d347, d348, d349, d350, d351, d352, d353, d354, d355, d356, d357, d358, d359, d360, d361, d362, d363, d364, d365, d366, d367, d368, d369, d370, d371, d372, d373, d374, d375, d376, d377, d378, d379, d380, d381, d382, d383, d384, d385, d386, d387, d388, d389, d390, d391, d392, d393, d394, d395, d396, d397, d398, d399, d400, d401, d402, d403, d404, d405, d406, d407, d408, d409, d410, d411, d412, d413, d414;

	not (d1, x3);
	xor (d2, x2);
	xor (d3, x4);
	nand (d4, x2, x3);
	xor (d5, x0, x3);
	and (d6, x0, x5);
	nor (d7, x0, x1);
	or (d8, x3, x5);
	buf (d9, x4);
	xnor (d10, x3, x5);
	nand (d11, x0, x4);
	or (d12, x1, x5);
	not (d13, x1);
	not (d14, x2);
	xor (d15, x0, x5);
	buf (d16, x3);
	xor (d17, x1);
	xor (d18, x0, x4);
	not (d19, x4);
	buf (d20, x0);
	nand (d21, x2, x5);
	xor (d22, x0, x2);
	and (d23, x2, x4);
	and (d24, x0, x2);
	xnor (d25, x3);
	nor (d26, x0, x4);
	buf (d27, x2);
	or (d28, x4, x5);
	xor (d29, x1, x4);
	or (d30, x3, x5);
	nor (d31, x0, x5);
	or (d32, d2, d24);
	or (d33, d31);
	nand (d34, d8, d31);
	or (d35, d29, d30);
	and (d36, d13, d25);
	xor (d37, d14);
	or (d38, d4, d14);
	nor (d39, d22);
	not (d40, d30);
	xnor (d41, d4, d23);
	nand (d42, d8);
	or (d43, d7);
	not (d44, d22);
	xor (d45, d25, d29);
	buf (d46, d25);
	buf (d47, d23);
	nand (d48, d15, d24);
	buf (d49, d1);
	xnor (d50, d4, d25);
	xor (d51, d15, d19);
	and (d52, d20, d27);
	nand (d53, d9, d11);
	buf (d54, d28);
	nand (d55, d12, d21);
	buf (d56, d15);
	and (d57, d24, d27);
	and (d58, d5, d16);
	xnor (d59, d6, d19);
	not (d60, x0);
	xnor (d61, d11, d16);
	nand (d62, d22, d26);
	xor (d63, d18, d20);
	not (d64, d2);
	not (d65, d19);
	xnor (d66, d18, d25);
	xor (d67, d5, d19);
	xor (d68, d4, d16);
	or (d69, d6, d14);
	nor (d70, d18, d30);
	nor (d71, d1, d18);
	buf (d72, d20);
	or (d73, d11, d22);
	or (d74, d13, d22);
	nand (d75, d5, d12);
	not (d76, d14);
	nand (d77, d8, d29);
	and (d78, d19, d25);
	xor (d79, d2, d25);
	xor (d80, d14, d22);
	buf (d81, d8);
	xnor (d82, d5, d25);
	buf (d83, d7);
	nor (d84, d38, d40);
	buf (d85, d74);
	and (d86, d54, d62);
	xnor (d87, d40, d52);
	or (d88, d52, d66);
	not (d89, d62);
	and (d90, d43, d76);
	or (d91, d42, d73);
	xor (d92, d32, d43);
	nand (d93, d42, d73);
	xor (d94, d40, d54);
	not (d95, d37);
	and (d96, d40, d74);
	buf (d97, d50);
	xnor (d98, d40, d72);
	nor (d99, d43, d50);
	nand (d100, d40, d57);
	or (d101, d32, d42);
	nor (d102, d92, d97);
	xnor (d103, d91, d101);
	nand (d104, d95, d96);
	and (d105, d99);
	xor (d106, d86, d93);
	not (d107, d94);
	xnor (d108, d92, d99);
	buf (d109, d16);
	buf (d110, x1);
	not (d111, d59);
	not (d112, d21);
	and (d113, d95);
	nand (d114, d88, d97);
	xnor (d115, d96, d99);
	buf (d116, d40);
	nand (d117, d86, d93);
	buf (d118, d61);
	or (d119, d89, d100);
	and (d120, d87, d98);
	or (d121, d88, d89);
	xor (d122, d92, d99);
	nand (d123, d89, d95);
	xnor (d124, d97, d101);
	xor (d125, d87, d89);
	nor (d126, d84, d95);
	not (d127, d13);
	xnor (d128, d88, d97);
	not (d129, d42);
	buf (d130, d67);
	nand (d131, d95, d98);
	nor (d132, d95, d98);
	nor (d133, d99, d100);
	or (d134, d85, d90);
	and (d135, d84, d98);
	buf (d136, d19);
	not (d137, d66);
	and (d138, d93, d101);
	buf (d139, d88);
	xor (d140, d83, d98);
	not (d141, d87);
	xnor (d142, d87, d94);
	buf (d143, d6);
	nand (d144, d85, d89);
	nand (d145, d93, d94);
	nand (d146, d83, d87);
	and (d147, d83, d100);
	not (d148, d47);
	not (d149, x5);
	nor (d150, d104, d141);
	xnor (d151, d109, d136);
	nand (d152, d118, d128);
	nor (d153, d103, d109);
	not (d154, d40);
	buf (d155, d49);
	not (d156, d115);
	and (d157, d110, d137);
	xor (d158, d109);
	xor (d159, d123, d133);
	nand (d160, d116, d124);
	or (d161, d126, d144);
	not (d162, d103);
	and (d163, d120, d142);
	nor (d164, d129, d143);
	xor (d165, d104, d135);
	not (d166, d20);
	or (d167, d111, d114);
	nor (d168, d132, d144);
	not (d169, d56);
	and (d170, d114, d140);
	or (d171, d108, d113);
	buf (d172, d118);
	or (d173, d109, d136);
	xor (d174, d110, d122);
	nand (d175, d107, d124);
	and (d176, d134, d147);
	nand (d177, d134, d146);
	nand (d178, d132, d136);
	and (d179, d120, d135);
	and (d180, d115, d133);
	and (d181, d105, d108);
	not (d182, d81);
	or (d183, d116, d123);
	not (d184, d58);
	xor (d185, d116, d139);
	xor (d186, d107, d141);
	not (d187, d125);
	xnor (d188, d104, d120);
	not (d189, d74);
	or (d190, d129, d130);
	nand (d191, d127, d144);
	or (d192, d114, d120);
	xnor (d193, d119, d136);
	nand (d194, d131);
	xnor (d195, d107, d137);
	nor (d196, d126, d128);
	xor (d197, d119, d139);
	buf (d198, d48);
	nand (d199, d138, d140);
	buf (d200, d107);
	xor (d201, d105, d141);
	and (d202, d126, d147);
	xor (d203, d123, d140);
	xnor (d204, d113, d144);
	not (d205, d133);
	xor (d206, d106, d146);
	and (d207, d108, d122);
	and (d208, d119, d120);
	nor (d209, d120, d122);
	buf (d210, d111);
	and (d211, d103, d108);
	not (d212, d129);
	or (d213, d121, d136);
	nor (d214, d132, d140);
	and (d215, d113, d139);
	buf (d216, d99);
	xor (d217, d126, d136);
	nand (d218, d108, d145);
	or (d219, d106, d131);
	or (d220, d103, d117);
	nand (d221, d109, d122);
	buf (d222, d60);
	not (d223, d27);
	not (d224, d128);
	nand (d225, d113, d118);
	xnor (d226, d126, d130);
	xor (d227, d159, d199);
	nor (d228, d150, d177);
	or (d229, d165, d166);
	nand (d230, d149, d191);
	buf (d231, d81);
	nand (d232, d197, d204);
	or (d233, d165, d169);
	xnor (d234, d156, d226);
	buf (d235, d193);
	xnor (d236, d229, d235);
	or (d237, d234, d235);
	or (d238, d227, d233);
	nand (d239, d229, d231);
	xnor (d240, d232, d234);
	nand (d241, d228, d234);
	nand (d242, d227, d231);
	and (d243, d229, d233);
	not (d244, d5);
	buf (d245, d69);
	nand (d246, d227);
	nor (d247, d230, d232);
	or (d248, d230, d234);
	and (d249, d228, d229);
	or (d250, d231, d233);
	buf (d251, d109);
	nand (d252, d231, d234);
	xor (d253, d229, d231);
	xnor (d254, d231, d233);
	xor (d255, d229, d233);
	not (d256, d156);
	and (d257, d227, d232);
	not (d258, d181);
	buf (d259, d59);
	xor (d260, d227, d235);
	xor (d261, d227, d234);
	not (d262, d121);
	xor (d263, d233, d235);
	nor (d264, d230, d233);
	buf (d265, d234);
	not (d266, d147);
	not (d267, d104);
	or (d268, d229, d234);
	and (d269, d232, d235);
	not (d270, d220);
	xnor (d271, d228, d230);
	nor (d272, d230, d235);
	xnor (d273, d230);
	nand (d274, d235);
	and (d275, d231, d235);
	xnor (d276, d244, d249);
	buf (d277, d161);
	nor (d278, d268, d274);
	or (d279, d239, d245);
	or (d280, d253, d264);
	nor (d281, d238, d275);
	xnor (d282, d255, d275);
	xnor (d283, d239, d264);
	buf (d284, d199);
	or (d285, d244, d265);
	xnor (d286, d262, d270);
	xor (d287, d241, d272);
	nor (d288, d251, d253);
	and (d289, d236, d263);
	and (d290, d236, d242);
	nand (d291, d240, d242);
	nor (d292, d237, d274);
	xnor (d293, d251, d255);
	xnor (d294, d256, d275);
	and (d295, d243, d271);
	buf (d296, d85);
	xor (d297, d267, d275);
	xnor (d298, d264, d269);
	not (d299, d109);
	buf (d300, d247);
	not (d301, d274);
	not (d302, d7);
	xnor (d303, d241, d265);
	buf (d304, d12);
	and (d305, d250, d252);
	xnor (d306, d240, d274);
	xnor (d307, d249, d273);
	nor (d308, d253);
	xnor (d309, d245, d274);
	nand (d310, d240, d243);
	nor (d311, d237, d245);
	and (d312, d236, d250);
	buf (d313, d130);
	or (d314, d246, d251);
	or (d315, d251, d253);
	nor (d316, d249, d268);
	and (d317, d247, d249);
	nand (d318, d236, d251);
	and (d319, d252, d267);
	and (d320, d243, d253);
	nand (d321, d250, d266);
	or (d322, d255, d274);
	xnor (d323, d244, d248);
	and (d324, d236, d237);
	buf (d325, d140);
	and (d326, d255, d262);
	nand (d327, d240, d247);
	nand (d328, d273);
	and (d329, d252, d260);
	nand (d330, d260, d267);
	xnor (d331, d270, d271);
	or (d332, d236, d262);
	and (d333, d267, d271);
	nand (d334, d262, d266);
	buf (d335, d37);
	nor (d336, d238, d267);
	xor (d337, d265, d269);
	nor (d338, d252, d269);
	or (d339, d245, d272);
	buf (d340, d166);
	buf (d341, d220);
	and (d342, d254, d266);
	not (d343, d210);
	nand (d344, d265, d274);
	nor (d345, d238, d273);
	nor (d346, d239, d253);
	and (d347, d248, d253);
	and (d348, d257, d259);
	and (d349, d242, d256);
	nand (d350, d265, d266);
	or (d351, d239, d245);
	and (d352, d298, d340);
	xor (d353, d292, d347);
	and (d354, d315, d336);
	not (d355, d186);
	or (d356, d294, d307);
	xnor (d357, d313, d341);
	xor (d358, d316, d335);
	nor (d359, d321, d322);
	or (d360, d344, d349);
	and (d361, d278, d302);
	and (d362, d277, d341);
	xor (d363, d306, d338);
	nand (d364, d290, d316);
	and (d365, d308, d349);
	buf (d366, d125);
	xor (d367, d297, d298);
	nand (d368, d303, d351);
	nand (d369, d299, d332);
	nand (d370, d310, d336);
	buf (d371, d86);
	not (d372, d9);
	xor (d373, d316, d338);
	xnor (d374, d301, d345);
	nor (d375, d328, d344);
	or (d376, d308, d348);
	nand (d377, d276, d335);
	nor (d378, d278, d293);
	and (d379, d309, d341);
	and (d380, d301, d339);
	xor (d381, d294, d312);
	nand (d382, d323, d329);
	nor (d383, d281, d309);
	and (d384, d341, d349);
	not (d385, d332);
	not (d386, d291);
	nand (d387, d327, d345);
	nor (d388, d302, d308);
	not (d389, d241);
	or (d390, d285, d335);
	and (d391, d297, d305);
	not (d392, d256);
	and (d393, d316, d329);
	nand (d394, d286, d348);
	xnor (d395, d281, d305);
	buf (d396, d13);
	buf (d397, d4);
	or (d398, d286, d307);
	or (d399, d310, d347);
	xor (d400, d290, d343);
	or (d401, d311, d312);
	xor (d402, d283, d291);
	nand (d403, d294, d331);
	xnor (d404, d283, d323);
	xor (d405, d329, d334);
	nor (d406, d286, d343);
	xnor (d407, d300, d315);
	or (d408, d280, d346);
	nand (d409, d281, d301);
	buf (d410, d250);
	nor (d411, d279, d317);
	buf (d412, d265);
	and (d413, d307, d343);
	buf (d414, d141);
	assign f1 = d390;
	assign f2 = d371;
	assign f3 = d372;
	assign f4 = d355;
	assign f5 = d395;
	assign f6 = d403;
	assign f7 = d392;
	assign f8 = d384;
	assign f9 = d373;
	assign f10 = d411;
	assign f11 = d386;
	assign f12 = d379;
	assign f13 = d406;
	assign f14 = d394;
endmodule
