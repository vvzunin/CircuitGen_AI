module CCGRCG34( x0, x1, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17, f18, f19 );

	input x0, x1;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17, f18, f19;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314, d315, d316, d317, d318, d319, d320, d321, d322, d323, d324, d325, d326, d327, d328, d329, d330, d331, d332, d333, d334, d335, d336, d337, d338, d339, d340, d341, d342, d343, d344, d345, d346, d347, d348, d349, d350, d351, d352, d353, d354, d355, d356, d357, d358, d359, d360, d361, d362, d363, d364, d365, d366, d367, d368, d369, d370, d371, d372, d373, d374, d375;

	xnor (d1, x0, x1);
	and (d2, x0);
	nor (d3, x0);
	xor (d4, x0);
	buf (d5, x0);
	buf (d6, x1);
	nor (d7, x0, x1);
	and (d8, x1);
	and (d9, x0, x1);
	not (d10, x1);
	nand (d11, x1);
	xnor (d12, x1);
	or (d13, x0, x1);
	or (d14, x0);
	xor (d15, x1);
	or (d16, x1);
	xor (d17, x0, x1);
	nor (d18, x1);
	and (d19, x0, x1);
	not (d20, x0);
	xnor (d21, x0);
	nand (d22, x0, x1);
	nor (d23, x0, x1);
	xor (d24, x0, x1);
	nand (d25, x0);
	or (d26, x0, x1);
	nand (d27, x0, x1);
	not (d28, d7);
	xnor (d29, d3, d12);
	xnor (d30, d11, d16);
	or (d31, d13, d14);
	or (d32, d23, d25);
	or (d33, d20, d25);
	xor (d34, d5, d25);
	nor (d35, d20);
	or (d36, d7, d19);
	or (d37, d7, d25);
	buf (d38, d7);
	xor (d39, d12, d26);
	xor (d40, d23, d27);
	buf (d41, d1);
	and (d42, d6, d23);
	xor (d43, d3, d11);
	buf (d44, d9);
	xor (d45, d12, d15);
	xnor (d46, d14, d16);
	nor (d47, d12, d15);
	or (d48, d5, d25);
	nand (d49, d14, d17);
	or (d50, d14, d25);
	xor (d51, d22, d23);
	nand (d52, d18, d23);
	or (d53, d18, d20);
	xor (d54, d22, d24);
	nor (d55, d13, d18);
	buf (d56, d3);
	not (d57, d5);
	buf (d58, d2);
	nand (d59, d18, d26);
	nor (d60, d7, d24);
	or (d61, d2, d19);
	xor (d62, d18, d20);
	or (d63, d1, d13);
	nor (d64, d5);
	and (d65, d2, d27);
	buf (d66, d14);
	nor (d67, d2, d26);
	nand (d68, d23);
	nand (d69, d16);
	xnor (d70, d3, d7);
	not (d71, d12);
	or (d72, d4, d10);
	nor (d73, d19, d26);
	nand (d74, d15, d16);
	nand (d75, d20, d21);
	buf (d76, d24);
	nand (d77, d11, d26);
	nor (d78, d10, d16);
	and (d79, d15, d26);
	xor (d80, d3, d22);
	xor (d81, d11, d19);
	or (d82, d16, d21);
	nand (d83, d4, d5);
	buf (d84, d23);
	or (d85, d24, d25);
	nor (d86, d1, d11);
	buf (d87, d22);
	nand (d88, d15, d27);
	xor (d89, d13, d26);
	not (d90, d8);
	not (d91, d18);
	buf (d92, d11);
	and (d93, d19, d22);
	and (d94, d1, d24);
	nor (d95, d8, d24);
	or (d96, d10, d23);
	nand (d97, d14, d20);
	xor (d98, d15, d27);
	buf (d99, d8);
	xnor (d100, d1, d21);
	and (d101, d9, d10);
	nor (d102, d10, d18);
	nor (d103, d14, d24);
	not (d104, d21);
	nor (d105, d15, d16);
	nor (d106, d23, d26);
	xor (d107, d39, d91);
	nand (d108, d29, d54);
	xor (d109, d29, d48);
	nand (d110, d84, d91);
	xnor (d111, d61, d92);
	buf (d112, d41);
	not (d113, d10);
	nor (d114, d68, d70);
	and (d115, d57, d58);
	xnor (d116, d36, d51);
	xnor (d117, d95, d97);
	or (d118, d70, d104);
	buf (d119, d39);
	xor (d120, d32, d76);
	nand (d121, d70, d106);
	nand (d122, d35, d49);
	not (d123, d34);
	xor (d124, d60, d73);
	or (d125, d45, d83);
	not (d126, d46);
	nand (d127, d42, d65);
	or (d128, d53, d92);
	and (d129, d32, d77);
	xnor (d130, d40, d58);
	not (d131, d84);
	xnor (d132, d92, d100);
	or (d133, d31, d45);
	xor (d134, d51, d97);
	nand (d135, d45, d103);
	xnor (d136, d87, d104);
	xor (d137, d54, d96);
	not (d138, d20);
	xnor (d139, d46, d74);
	and (d140, d41, d81);
	nand (d141, d103, d104);
	xor (d142, d45, d48);
	xor (d143, d71, d80);
	xor (d144, d36, d44);
	not (d145, d13);
	xnor (d146, d46, d57);
	nand (d147, d57, d91);
	nor (d148, d37, d65);
	xor (d149, d41, d75);
	buf (d150, d20);
	or (d151, d58, d90);
	or (d152, d56, d57);
	nor (d153, d43, d78);
	xnor (d154, d61, d62);
	nor (d155, d44, d71);
	nand (d156, d44, d70);
	or (d157, d50, d69);
	not (d158, d79);
	not (d159, d95);
	xor (d160, d55, d77);
	buf (d161, d74);
	nor (d162, d47, d70);
	buf (d163, d44);
	xnor (d164, d49, d87);
	nor (d165, d30, d67);
	nor (d166, d31, d53);
	buf (d167, d90);
	xnor (d168, d38, d66);
	xnor (d169, d55, d84);
	xnor (d170, d64, d73);
	xor (d171, d60, d97);
	xnor (d172, d80, d82);
	or (d173, d65, d96);
	or (d174, d95, d102);
	and (d175, d34, d74);
	or (d176, d43, d79);
	buf (d177, d54);
	nand (d178, d28, d99);
	nor (d179, d29, d81);
	not (d180, d53);
	buf (d181, d6);
	nand (d182, d36, d87);
	nand (d183, d53, d92);
	xor (d184, d50, d89);
	xnor (d185, d38, d96);
	xor (d186, d82, d87);
	and (d187, d43, d94);
	and (d188, d62, d91);
	xnor (d189, d35, d105);
	or (d190, d47, d80);
	xor (d191, d76, d89);
	nand (d192, d28, d105);
	xor (d193, d31, d94);
	xor (d194, d80, d101);
	not (d195, d66);
	xor (d196, d156, d177);
	nor (d197, d120, d181);
	not (d198, d97);
	xnor (d199, d155, d182);
	xor (d200, d120, d144);
	not (d201, d36);
	xor (d202, d169, d191);
	or (d203, d134, d185);
	and (d204, d148, d166);
	not (d205, d161);
	xnor (d206, d138, d190);
	nand (d207, d109, d159);
	and (d208, d145, d155);
	nand (d209, d174, d177);
	nor (d210, d114, d145);
	and (d211, d171, d179);
	xor (d212, d108, d123);
	or (d213, d157, d166);
	xor (d214, d122, d127);
	or (d215, d115, d164);
	xor (d216, d114, d184);
	or (d217, d133, d187);
	or (d218, d171, d191);
	not (d219, d153);
	xnor (d220, d129, d166);
	xnor (d221, d118, d181);
	xnor (d222, d145, d190);
	and (d223, d111, d190);
	and (d224, d162, d175);
	nor (d225, d138, d166);
	not (d226, d23);
	or (d227, d152, d163);
	buf (d228, d188);
	and (d229, d173, d184);
	buf (d230, d190);
	xor (d231, d170, d173);
	buf (d232, d116);
	nand (d233, d152, d169);
	xnor (d234, d143, d163);
	and (d235, d126, d183);
	not (d236, d160);
	xnor (d237, d114, d132);
	nand (d238, d129, d161);
	or (d239, d132, d156);
	xor (d240, d122, d163);
	xor (d241, d130, d159);
	not (d242, d81);
	xnor (d243, d108, d164);
	xnor (d244, d149, d165);
	nand (d245, d138, d173);
	and (d246, d117, d185);
	xnor (d247, d168, d181);
	nand (d248, d137, d173);
	and (d249, d172, d190);
	xor (d250, d151, d154);
	xor (d251, d132, d142);
	buf (d252, d185);
	buf (d253, d121);
	or (d254, d121, d183);
	buf (d255, d31);
	xnor (d256, d177, d194);
	buf (d257, d95);
	xnor (d258, d148, d187);
	xnor (d259, d199, d230);
	not (d260, d231);
	not (d261, d96);
	not (d262, d223);
	nand (d263, d198, d218);
	or (d264, d238, d240);
	or (d265, d223, d255);
	or (d266, d206, d235);
	nor (d267, d207, d253);
	nor (d268, d205, d220);
	nand (d269, d200, d205);
	not (d270, d99);
	xor (d271, d229, d241);
	or (d272, d204, d213);
	not (d273, d217);
	nor (d274, d199, d225);
	and (d275, d221, d231);
	and (d276, d210, d254);
	or (d277, d206, d221);
	and (d278, d204, d217);
	xor (d279, d224, d256);
	and (d280, d196, d233);
	or (d281, d242, d251);
	xor (d282, d219, d253);
	not (d283, d51);
	nand (d284, d201, d236);
	xnor (d285, d201, d221);
	and (d286, d198, d219);
	nand (d287, d197, d217);
	buf (d288, d241);
	nand (d289, d230, d247);
	xnor (d290, d197, d201);
	buf (d291, d124);
	nand (d292, d218, d250);
	buf (d293, d62);
	not (d294, d48);
	nand (d295, d203, d240);
	not (d296, d172);
	not (d297, d37);
	xor (d298, d225, d242);
	or (d299, d204, d215);
	nor (d300, d204, d226);
	not (d301, d9);
	and (d302, d210, d232);
	or (d303, d224, d230);
	nor (d304, d227, d251);
	nand (d305, d236, d248);
	xnor (d306, d208, d224);
	nor (d307, d225, d234);
	and (d308, d248, d252);
	not (d309, d162);
	and (d310, d203, d204);
	buf (d311, d183);
	nor (d312, d248, d251);
	nand (d313, d197, d258);
	xor (d314, d235, d256);
	xor (d315, d222, d257);
	or (d316, d204, d219);
	buf (d317, d181);
	or (d318, d253);
	nor (d319, d250, d256);
	nor (d320, d236, d249);
	xnor (d321, d201, d232);
	xor (d322, d264, d273);
	not (d323, d265);
	or (d324, d305, d314);
	and (d325, d319, d321);
	or (d326, d314, d316);
	buf (d327, d46);
	buf (d328, d282);
	xnor (d329, d276, d282);
	or (d330, d260, d309);
	xor (d331, d282, d285);
	or (d332, d273, d301);
	not (d333, d38);
	buf (d334, d162);
	nand (d335, d277, d316);
	or (d336, d267, d315);
	xnor (d337, d259, d282);
	or (d338, d271, d286);
	buf (d339, d257);
	nand (d340, d295, d308);
	and (d341, d317, d321);
	not (d342, d244);
	or (d343, d299, d319);
	nand (d344, d295, d302);
	and (d345, d281, d316);
	or (d346, d296, d315);
	nand (d347, d266, d267);
	and (d348, d281, d285);
	or (d349, d276, d283);
	or (d350, d318, d321);
	xnor (d351, d307, d315);
	xor (d352, d263, d309);
	buf (d353, d269);
	nor (d354, d278, d290);
	buf (d355, d77);
	or (d356, d298, d318);
	not (d357, d284);
	xor (d358, d284, d315);
	not (d359, d43);
	xnor (d360, d290, d316);
	xor (d361, d315, d321);
	or (d362, d298, d318);
	and (d363, d286, d296);
	and (d364, d288, d295);
	xnor (d365, d302, d305);
	or (d366, d278, d305);
	xnor (d367, d277, d304);
	buf (d368, d199);
	nand (d369, d266, d291);
	xnor (d370, d260, d286);
	xnor (d371, d268, d321);
	xnor (d372, d274, d275);
	and (d373, d276, d296);
	nand (d374, d311, d317);
	nor (d375, d272, d284);
	assign f1 = d322;
	assign f2 = d363;
	assign f3 = d347;
	assign f4 = d364;
	assign f5 = d360;
	assign f6 = d359;
	assign f7 = d367;
	assign f8 = d346;
	assign f9 = d337;
	assign f10 = d330;
	assign f11 = d366;
	assign f12 = d347;
	assign f13 = d357;
	assign f14 = d374;
	assign f15 = d347;
	assign f16 = d348;
	assign f17 = d347;
	assign f18 = d326;
	assign f19 = d341;
endmodule
