module CCGRCG20( x0, x1, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12 );

	input x0, x1;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314, d315, d316, d317, d318, d319, d320, d321, d322, d323, d324, d325, d326, d327, d328, d329, d330, d331, d332, d333, d334, d335, d336, d337, d338, d339, d340;

	or (d1, x1);
	nor (d2, x1);
	buf (d3, x1);
	or (d4, x0, x1);
	nand (d5, x0, x1);
	and (d6, x0);
	not (d7, x0);
	xnor (d8, x0, x1);
	xor (d9, x0);
	not (d10, x1);
	and (d11, x1);
	or (d12, x0, x1);
	and (d13, x0, x1);
	nor (d14, x0, x1);
	xor (d15, x0, x1);
	xnor (d16, x0);
	nand (d17, x0);
	xnor (d18, x0, x1);
	xor (d19, x0, x1);
	xnor (d20, x1);
	buf (d21, x0);
	xor (d22, x1);
	or (d23, d19, d20);
	xor (d24, d2, d4);
	or (d25, d3, d10);
	not (d26, d9);
	nand (d27, d5, d19);
	nand (d28, d1, d3);
	or (d29, d4, d18);
	nor (d30, d4, d17);
	nor (d31, d20, d22);
	and (d32, d2, d18);
	xor (d33, d9, d10);
	xor (d34, d1, d13);
	xnor (d35, d1, d11);
	or (d36, d6, d12);
	xor (d37, d8, d18);
	xor (d38, d18, d19);
	nand (d39, d15, d16);
	xnor (d40, d6, d15);
	not (d41, d17);
	and (d42, d25, d36);
	or (d43, d24, d38);
	xor (d44, d23, d34);
	nand (d45, d39, d40);
	xor (d46, d24, d30);
	xor (d47, d28, d39);
	buf (d48, d40);
	or (d49, d25, d32);
	buf (d50, d22);
	nand (d51, d23, d32);
	and (d52, d23, d28);
	or (d53, d31, d33);
	buf (d54, d6);
	or (d55, d24, d29);
	xor (d56, d28, d40);
	nor (d57, d23, d40);
	or (d58, d28, d31);
	and (d59, d25, d28);
	and (d60, d27, d33);
	or (d61, d28, d34);
	or (d62, d24, d39);
	buf (d63, d23);
	xor (d64, d32, d34);
	xor (d65, d32, d35);
	and (d66, d30, d39);
	xnor (d67, d28, d40);
	nor (d68, d26, d32);
	xor (d69, d32, d38);
	xor (d70, d24, d26);
	buf (d71, d13);
	not (d72, d2);
	or (d73, d31, d32);
	nor (d74, d29, d36);
	xor (d75, d36);
	nand (d76, d25, d33);
	not (d77, d7);
	nand (d78, d23);
	not (d79, d36);
	buf (d80, d17);
	buf (d81, d3);
	and (d82, d26, d34);
	and (d83, d30, d34);
	nor (d84, d40);
	xor (d85, d30, d40);
	xnor (d86, d24, d38);
	buf (d87, d2);
	xnor (d88, d31, d33);
	and (d89, d36, d37);
	nor (d90, d26, d40);
	nand (d91, d24, d39);
	and (d92, d27, d37);
	buf (d93, d28);
	buf (d94, d34);
	xnor (d95, d32, d35);
	nand (d96, d29, d38);
	and (d97, d26, d29);
	nor (d98, d30, d38);
	xnor (d99, d31, d39);
	xnor (d100, d31, d38);
	buf (d101, d12);
	nor (d102, d27, d30);
	nor (d103, d38);
	or (d104, d30, d37);
	nand (d105, d31, d40);
	xnor (d106, d33, d38);
	xnor (d107, d32, d40);
	not (d108, d4);
	and (d109, d25, d36);
	and (d110, d29, d32);
	nand (d111, d26, d36);
	and (d112, d32);
	buf (d113, d8);
	xor (d114, d32, d40);
	xnor (d115, d26, d34);
	nand (d116, d23, d35);
	xnor (d117, d38);
	or (d118, d28, d33);
	and (d119, d33, d39);
	xor (d120, d30, d33);
	nand (d121, d53, d90);
	nand (d122, d44, d49);
	xor (d123, d93, d111);
	nand (d124, d66, d89);
	and (d125, d72, d94);
	xnor (d126, d91, d95);
	not (d127, d84);
	nor (d128, d71, d97);
	not (d129, d37);
	buf (d130, d97);
	buf (d131, d99);
	buf (d132, d58);
	nand (d133, d72, d117);
	xnor (d134, d58, d120);
	nand (d135, d54, d84);
	nand (d136, d41, d66);
	nand (d137, d76, d118);
	or (d138, d42, d79);
	or (d139, d129, d133);
	not (d140, d100);
	nor (d141, d130, d136);
	or (d142, d121, d125);
	xnor (d143, d126, d131);
	nand (d144, d131, d137);
	not (d145, d72);
	not (d146, d110);
	xor (d147, d133, d134);
	nand (d148, d133, d135);
	not (d149, d54);
	not (d150, d31);
	not (d151, d81);
	buf (d152, d88);
	and (d153, d128, d137);
	xor (d154, d123, d133);
	nor (d155, d130, d138);
	xor (d156, d123, d134);
	xnor (d157, d125, d127);
	buf (d158, d26);
	nor (d159, d132, d133);
	buf (d160, d33);
	xnor (d161, d125, d126);
	nand (d162, d123, d125);
	nor (d163, d129, d136);
	not (d164, d85);
	or (d165, d121, d134);
	and (d166, d126, d133);
	not (d167, d79);
	and (d168, d122, d133);
	or (d169, d126, d132);
	not (d170, d70);
	xor (d171, d125, d135);
	xor (d172, d134, d136);
	xnor (d173, d123, d135);
	buf (d174, d132);
	nor (d175, d130, d131);
	nand (d176, d122, d138);
	xnor (d177, d124, d130);
	xor (d178, d124, d134);
	xor (d179, d127, d135);
	xnor (d180, d131, d135);
	not (d181, d103);
	xnor (d182, d127, d138);
	xnor (d183, d126, d130);
	and (d184, d129, d131);
	nand (d185, d129, d137);
	and (d186, d123, d126);
	nand (d187, d130, d134);
	nor (d188, d128, d138);
	and (d189, d129, d131);
	and (d190, d125, d138);
	and (d191, d128, d132);
	and (d192, d122, d129);
	buf (d193, d53);
	nand (d194, d121, d138);
	buf (d195, d91);
	or (d196, d125, d126);
	or (d197, d133, d136);
	or (d198, d123, d135);
	not (d199, d89);
	and (d200, d125, d130);
	not (d201, d130);
	xnor (d202, d129, d138);
	nand (d203, d132, d137);
	and (d204, d123, d133);
	or (d205, d129, d132);
	nand (d206, d122, d134);
	xnor (d207, d134, d136);
	nand (d208, d122, d138);
	or (d209, d122, d135);
	nor (d210, d125, d132);
	or (d211, d125, d137);
	or (d212, d124, d131);
	not (d213, d90);
	nor (d214, d131, d137);
	buf (d215, d15);
	and (d216, d182, d188);
	buf (d217, d183);
	not (d218, d118);
	xor (d219, d154, d155);
	nand (d220, d152, d173);
	xnor (d221, d186, d198);
	not (d222, d167);
	buf (d223, d180);
	xnor (d224, d196, d201);
	xnor (d225, d162, d184);
	nor (d226, d154, d173);
	nand (d227, d163, d186);
	not (d228, d137);
	and (d229, d172, d210);
	xor (d230, d166, d210);
	nand (d231, d152, d190);
	xnor (d232, d153, d157);
	or (d233, d167, d177);
	nor (d234, d159, d161);
	xnor (d235, d160);
	or (d236, d180, d207);
	xor (d237, d168, d185);
	xor (d238, d160, d163);
	xnor (d239, d163, d171);
	nor (d240, d158, d187);
	xnor (d241, d162, d164);
	nand (d242, d153, d199);
	nor (d243, d147, d178);
	or (d244, d143, d178);
	xnor (d245, d148, d171);
	and (d246, d151, d179);
	nand (d247, d149, d193);
	xnor (d248, d144, d188);
	and (d249, d182, d194);
	or (d250, d147, d154);
	not (d251, d29);
	or (d252, d180, d211);
	nand (d253, d172, d212);
	nor (d254, d181, d196);
	nor (d255, d225, d230);
	xor (d256, d225, d254);
	xor (d257, d230, d243);
	xor (d258, d231, d245);
	and (d259, d229, d237);
	xnor (d260, d238, d252);
	and (d261, d229, d252);
	buf (d262, d18);
	and (d263, d222, d231);
	buf (d264, d187);
	buf (d265, d191);
	xor (d266, d224, d248);
	nor (d267, d235, d249);
	and (d268, d224, d231);
	xor (d269, d232, d233);
	xnor (d270, d219, d246);
	and (d271, d230, d239);
	not (d272, d61);
	buf (d273, d254);
	nand (d274, d241, d248);
	buf (d275, d249);
	nand (d276, d237, d251);
	not (d277, d217);
	not (d278, d233);
	and (d279, d220, d221);
	buf (d280, d43);
	xor (d281, d220, d228);
	xor (d282, d227, d235);
	nand (d283, d217, d223);
	nor (d284, d229, d237);
	and (d285, d220, d245);
	or (d286, d220, d249);
	not (d287, d105);
	xnor (d288, d222, d238);
	nand (d289, d222, d242);
	xnor (d290, d232, d246);
	buf (d291, d126);
	or (d292, d237, d249);
	nand (d293, d227, d236);
	buf (d294, d39);
	xnor (d295, d235, d237);
	not (d296, d198);
	or (d297, d240, d248);
	and (d298, d242, d244);
	xnor (d299, d238, d245);
	and (d300, d219, d231);
	xnor (d301, d220, d235);
	or (d302, d234, d245);
	xor (d303, d228, d253);
	xnor (d304, d223, d248);
	or (d305, d220, d222);
	nand (d306, d217, d219);
	or (d307, d230, d254);
	not (d308, d25);
	or (d309, d220, d231);
	or (d310, d223, d234);
	xnor (d311, d229, d245);
	xor (d312, d216, d238);
	and (d313, d216, d241);
	nand (d314, d231, d234);
	not (d315, d190);
	xnor (d316, d241, d242);
	xor (d317, d216, d221);
	not (d318, d126);
	xor (d319, d223, d252);
	xnor (d320, d223, d241);
	nor (d321, d231, d240);
	xor (d322, d221, d231);
	not (d323, d152);
	xnor (d324, d254);
	and (d325, d230, d245);
	not (d326, d213);
	and (d327, d222, d252);
	nand (d328, d242, d244);
	xor (d329, d230, d245);
	nor (d330, d222, d234);
	buf (d331, d46);
	and (d332, d237, d253);
	and (d333, d245, d249);
	and (d334, d240, d244);
	or (d335, d230, d242);
	or (d336, d218, d232);
	nor (d337, d245, d251);
	buf (d338, d251);
	xor (d339, d238, d254);
	xnor (d340, d219, d225);
	assign f1 = d326;
	assign f2 = d259;
	assign f3 = d319;
	assign f4 = d281;
	assign f5 = d327;
	assign f6 = d325;
	assign f7 = d255;
	assign f8 = d332;
	assign f9 = d256;
	assign f10 = d281;
	assign f11 = d265;
	assign f12 = d332;
endmodule
