module CCGRCG88( x0, x1, x2, x3, f1, f2, f3, f4, f5, f6, f7, f8 );

	input x0, x1, x2, x3;
	output f1, f2, f3, f4, f5, f6, f7, f8;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92;

	nand (d1, x0, x2);
	or (d2, x1, x3);
	not (d3, x2);
	xor (d4, x0, x1);
	and (d5, x2, x3);
	not (d6, x3);
	nor (d7, x2, x3);
	and (d8, x0, x1);
	nand (d9, x0, x2);
	or (d10, x1, x2);
	xor (d11, x0, x1);
	buf (d12, x3);
	and (d13, x1, x2);
	buf (d14, x1);
	nand (d15, x1, x3);
	not (d16, d2);
	and (d17, d4, d7);
	xnor (d18, d5, d8);
	xor (d19, d11);
	not (d20, d8);
	or (d21, d1, d6);
	xor (d22, d2, d10);
	or (d23, d12, d14);
	buf (d24, x0);
	nor (d25, d2, d4);
	and (d26, d9, d10);
	or (d27, d4, d13);
	nor (d28, d5, d12);
	or (d29, d4, d5);
	xnor (d30, d6, d9);
	or (d31, d11, d15);
	xnor (d32, d2, d7);
	xor (d33, d10, d12);
	not (d34, d5);
	or (d35, d5, d10);
	nor (d36, d2, d15);
	nor (d37, d2, d5);
	nor (d38, d5, d12);
	and (d39, d2, d15);
	or (d40, d2, d14);
	and (d41, d3, d4);
	nand (d42, d1, d14);
	xnor (d43, d5, d6);
	and (d44, d33, d42);
	and (d45, d20, d38);
	buf (d46, d19);
	nor (d47, d19, d39);
	xnor (d48, d16, d39);
	nor (d49, d39, d42);
	nand (d50, d28, d39);
	nor (d51, d39, d43);
	not (d52, d17);
	xnor (d53, d24, d39);
	and (d54, d20, d30);
	and (d55, d24, d33);
	or (d56, d34, d38);
	or (d57, d26, d37);
	buf (d58, d2);
	xnor (d59, d28, d43);
	buf (d60, d5);
	and (d61, d18, d29);
	xor (d62, d32);
	xor (d63, d24, d29);
	xnor (d64, d27, d29);
	xor (d65, d30, d43);
	nor (d66, d32, d34);
	nand (d67, d23, d24);
	xnor (d68, d31, d40);
	not (d69, d18);
	nor (d70, d38);
	xnor (d71, d30, d38);
	nand (d72, d22, d33);
	nand (d73, d23, d31);
	nor (d74, d32, d34);
	nor (d75, d20);
	and (d76, d19, d42);
	not (d77, d37);
	buf (d78, d42);
	not (d79, d16);
	nand (d80, d19, d35);
	xor (d81, d16, d28);
	xnor (d82, d32, d43);
	nor (d83, d21, d37);
	and (d84, d19, d31);
	xor (d85, d19, d27);
	buf (d86, d29);
	not (d87, d7);
	nor (d88, d31, d34);
	not (d89, d31);
	xnor (d90, d18, d25);
	and (d91, d18, d33);
	buf (d92, d11);
	assign f1 = d51;
	assign f2 = d46;
	assign f3 = d77;
	assign f4 = d80;
	assign f5 = d53;
	assign f6 = d54;
	assign f7 = d60;
	assign f8 = d49;
endmodule
