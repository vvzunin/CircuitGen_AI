module CCGRCG118( x0, x1, x2, x3, x4, f1, f2, f3, f4 );

	input x0, x1, x2, x3, x4;
	output f1, f2, f3, f4;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314, d315, d316, d317, d318, d319, d320, d321, d322, d323, d324, d325, d326, d327, d328, d329, d330, d331, d332, d333, d334, d335, d336, d337, d338, d339, d340, d341, d342, d343, d344, d345, d346, d347, d348, d349, d350, d351, d352, d353, d354, d355, d356, d357, d358, d359, d360, d361, d362, d363, d364, d365, d366, d367, d368, d369, d370, d371, d372, d373, d374, d375, d376, d377, d378, d379, d380, d381, d382, d383, d384, d385, d386, d387, d388, d389, d390, d391, d392, d393, d394, d395, d396, d397, d398, d399, d400, d401, d402, d403, d404, d405, d406, d407, d408, d409, d410, d411, d412, d413, d414, d415, d416, d417, d418, d419;

	xnor (d1, x2, x4);
	nor (d2, x0);
	or (d3, x1, x4);
	nor (d4, x0, x4);
	or (d5, x1, x4);
	nand (d6, x0, x2);
	and (d7, x3, x4);
	nor (d8, x0, x1);
	not (d9, x0);
	or (d10, x0, x1);
	and (d11, x0, x4);
	nand (d12, x2, x3);
	or (d13, x3, x4);
	not (d14, x4);
	nand (d15, x0, x1);
	and (d16, x1, x2);
	and (d17, x0, x3);
	nand (d18, x1, x3);
	xor (d19, x1, x2);
	nor (d20, x1, x4);
	nand (d21, x0, x4);
	xor (d22, x0, x3);
	xnor (d23, x0, x2);
	nor (d24, x2, x3);
	xor (d25, x1, x4);
	nand (d26, x1);
	buf (d27, x2);
	or (d28, x2, x3);
	or (d29, x2, x4);
	and (d30, x1);
	buf (d31, x0);
	nand (d32, x1, x2);
	nand (d33, x0, x2);
	and (d34, x4);
	and (d35, x0, x1);
	xnor (d36, x0);
	and (d37, x0, x1);
	xor (d38, x1, x2);
	nand (d39, x0);
	xnor (d40, x3);
	buf (d41, x3);
	or (d42, x0);
	nand (d43, x0, x1);
	not (d44, x2);
	xor (d45, x2, x4);
	nand (d46, x2, x4);
	xnor (d47, x3, x4);
	xor (d48, x0, x3);
	and (d49, x2, x4);
	and (d50, x0);
	xor (d51, x4);
	xnor (d52, x0, x2);
	not (d53, x1);
	and (d54, x3, x4);
	xnor (d55, x0, x4);
	and (d56, d18, d48);
	nand (d57, d31, d50);
	nand (d58, d9, d28);
	nor (d59, d32, d54);
	nand (d60, d31, d40);
	xnor (d61, d15, d41);
	nand (d62, d25, d37);
	nor (d63, d33, d55);
	xor (d64, d6, d27);
	xnor (d65, d31, d54);
	nor (d66, d27, d31);
	nor (d67, d7, d15);
	xor (d68, d6, d22);
	nor (d69, d3, d51);
	buf (d70, d31);
	and (d71, d8, d46);
	and (d72, d22, d29);
	nor (d73, d6, d9);
	or (d74, d21, d27);
	or (d75, d22, d53);
	or (d76, d12, d52);
	nand (d77, d4, d14);
	nor (d78, d26, d48);
	xor (d79, d47, d53);
	xnor (d80, d6, d19);
	xor (d81, d24, d39);
	xor (d82, d4, d15);
	xnor (d83, d60, d78);
	xnor (d84, d65, d80);
	nand (d85, d67, d76);
	xnor (d86, d74, d81);
	or (d87, d62, d77);
	xor (d88, d67, d76);
	not (d89, d78);
	nand (d90, d57, d76);
	nor (d91, d64, d66);
	and (d92, d68, d74);
	nand (d93, d61, d66);
	xor (d94, d71, d79);
	nand (d95, d69, d76);
	buf (d96, d79);
	and (d97, d56, d57);
	nor (d98, d75);
	or (d99, d63, d65);
	nand (d100, d65, d72);
	not (d101, d55);
	xor (d102, d76, d82);
	and (d103, d71, d79);
	and (d104, d73, d82);
	and (d105, d62, d66);
	nand (d106, d74, d78);
	or (d107, d63, d72);
	buf (d108, d6);
	buf (d109, d24);
	or (d110, d58, d65);
	nor (d111, d63, d67);
	nor (d112, d61, d78);
	nand (d113, d58, d79);
	or (d114, d58, d69);
	or (d115, d64, d79);
	xnor (d116, d59, d61);
	xor (d117, d60, d67);
	xor (d118, d70, d78);
	buf (d119, d20);
	nor (d120, d56, d63);
	xnor (d121, d62, d64);
	nand (d122, d60, d65);
	nor (d123, d57, d75);
	xor (d124, d58, d70);
	xor (d125, d65, d66);
	nor (d126, d64, d71);
	and (d127, d64, d76);
	nor (d128, d68, d82);
	nand (d129, d60, d80);
	not (d130, d29);
	xnor (d131, d65, d74);
	not (d132, d25);
	buf (d133, d58);
	nand (d134, d77, d79);
	nand (d135, d63, d71);
	or (d136, d60, d70);
	and (d137, d65, d78);
	not (d138, d15);
	not (d139, d80);
	nor (d140, d58, d74);
	nor (d141, d65, d72);
	or (d142, d60, d80);
	and (d143, d61, d71);
	nor (d144, d62, d81);
	not (d145, d14);
	buf (d146, d39);
	nor (d147, d74, d77);
	xor (d148, d58, d68);
	or (d149, d63, d78);
	and (d150, d56, d71);
	not (d151, d31);
	nor (d152, d66, d80);
	not (d153, d33);
	nand (d154, d62, d68);
	nor (d155, d97, d115);
	xnor (d156, d101, d132);
	xor (d157, d120, d132);
	xnor (d158, d105, d121);
	buf (d159, d153);
	and (d160, d88, d95);
	nor (d161, d118, d150);
	nor (d162, d95, d140);
	not (d163, d53);
	xnor (d164, d97, d136);
	and (d165, d89, d123);
	nand (d166, d101, d109);
	nand (d167, d117, d124);
	nor (d168, d115, d119);
	buf (d169, d116);
	nor (d170, d96, d116);
	nor (d171, d87, d129);
	nor (d172, d114, d129);
	nor (d173, d148, d153);
	not (d174, d38);
	nand (d175, d117, d125);
	or (d176, d109, d113);
	xnor (d177, d136, d144);
	or (d178, d114, d139);
	not (d179, d108);
	nand (d180, d135, d150);
	and (d181, d83, d106);
	or (d182, d83, d106);
	xnor (d183, d133, d149);
	xnor (d184, d98, d146);
	nand (d185, d84, d125);
	nand (d186, d133, d146);
	and (d187, d95, d109);
	xor (d188, d117, d124);
	nor (d189, d105, d143);
	or (d190, d87, d120);
	and (d191, d92, d114);
	nand (d192, d123, d125);
	xnor (d193, d135);
	and (d194, d95, d122);
	buf (d195, d90);
	nand (d196, d152, d153);
	nand (d197, d101, d148);
	or (d198, d119, d144);
	or (d199, d110, d150);
	buf (d200, d137);
	and (d201, d165, d184);
	xor (d202, d181, d186);
	and (d203, d160, d171);
	and (d204, d163, d170);
	or (d205, d161, d194);
	nand (d206, d160, d184);
	or (d207, d159, d185);
	xor (d208, d177, d183);
	not (d209, d32);
	xor (d210, d179, d194);
	nor (d211, d156, d182);
	nand (d212, d159, d161);
	xnor (d213, d160, d190);
	buf (d214, d14);
	not (d215, d195);
	nand (d216, d172, d183);
	xor (d217, d161, d179);
	nor (d218, d189, d193);
	xor (d219, d181);
	nand (d220, d158, d196);
	nand (d221, d165, d166);
	xor (d222, d179, d194);
	nor (d223, d166, d169);
	xor (d224, d188, d189);
	and (d225, d162, d197);
	and (d226, d163, d187);
	or (d227, d178, d183);
	buf (d228, d113);
	xor (d229, d180, d192);
	not (d230, d39);
	nand (d231, d187);
	xnor (d232, d166, d167);
	not (d233, d165);
	or (d234, d172, d173);
	and (d235, d162, d176);
	and (d236, d164, d176);
	not (d237, d148);
	nand (d238, d173, d180);
	nor (d239, d157, d171);
	and (d240, d166, d176);
	buf (d241, d121);
	xor (d242, d162, d169);
	not (d243, d50);
	xor (d244, d172, d187);
	buf (d245, d114);
	or (d246, d158, d187);
	xnor (d247, d165, d178);
	or (d248, d167, d188);
	nor (d249, d195, d198);
	nand (d250, d170, d181);
	and (d251, d170, d171);
	not (d252, d57);
	nand (d253, d156, d180);
	xnor (d254, d168, d196);
	xor (d255, d159, d183);
	or (d256, d160, d197);
	nor (d257, d157, d160);
	nor (d258, d167, d189);
	buf (d259, d148);
	or (d260, d158, d199);
	xor (d261, d186, d191);
	buf (d262, d160);
	nor (d263, d176, d193);
	and (d264, d192, d197);
	not (d265, d43);
	nand (d266, d223, d256);
	xor (d267, d204, d247);
	and (d268, d215, d236);
	nand (d269, d226, d246);
	and (d270, d227, d256);
	buf (d271, d189);
	or (d272, d211, d254);
	buf (d273, d199);
	or (d274, d207, d259);
	nor (d275, d234, d247);
	and (d276, d239, d255);
	not (d277, d202);
	nand (d278, d216, d232);
	nor (d279, d220, d235);
	nand (d280, d255, d261);
	and (d281, d225, d257);
	not (d282, d62);
	and (d283, d210, d250);
	xnor (d284, d247, d259);
	nor (d285, d205, d251);
	nand (d286, d256, d260);
	nor (d287, d218, d261);
	nand (d288, d215, d217);
	nand (d289, d203, d212);
	buf (d290, d225);
	nand (d291, d211, d225);
	xnor (d292, d216, d226);
	or (d293, d218, d227);
	xnor (d294, d208, d247);
	xnor (d295, d215, d221);
	xor (d296, d224, d257);
	nand (d297, d235, d252);
	xnor (d298, d222, d250);
	not (d299, d223);
	not (d300, d26);
	or (d301, d207, d253);
	not (d302, d184);
	nor (d303, d238);
	xnor (d304, d237, d254);
	and (d305, d230, d260);
	and (d306, d204, d214);
	not (d307, d190);
	nand (d308, d216, d225);
	xor (d309, d214, d232);
	xor (d310, d241, d242);
	or (d311, d229, d260);
	xnor (d312, d240, d264);
	nand (d313, d250, d258);
	xor (d314, d217, d258);
	xnor (d315, d208, d243);
	xor (d316, d226, d230);
	and (d317, d213, d234);
	nor (d318, d244, d250);
	nand (d319, d216, d234);
	xor (d320, d241, d249);
	xnor (d321, d213, d263);
	buf (d322, d38);
	nand (d323, d213, d258);
	xnor (d324, d225, d232);
	xnor (d325, d209, d250);
	xor (d326, d233, d239);
	nor (d327, d220, d245);
	xnor (d328, d206, d250);
	nand (d329, d220, d226);
	not (d330, d171);
	or (d331, d219, d260);
	nand (d332, d235, d238);
	not (d333, d106);
	nand (d334, d211, d258);
	or (d335, d206, d257);
	nor (d336, d247, d264);
	nor (d337, d245);
	nor (d338, d226, d229);
	xnor (d339, d211, d240);
	and (d340, d222, d247);
	and (d341, d226, d250);
	nand (d342, d235, d253);
	or (d343, d212, d244);
	nor (d344, d225);
	or (d345, d261, d265);
	buf (d346, d122);
	xnor (d347, d236, d256);
	or (d348, d221, d222);
	nand (d349, d237, d245);
	nor (d350, d203, d207);
	or (d351, d204, d234);
	xor (d352, d219, d236);
	nor (d353, d277, d280);
	buf (d354, d245);
	nand (d355, d315, d346);
	xnor (d356, d288, d334);
	xor (d357, d267, d271);
	and (d358, d310, d344);
	xnor (d359, d293, d341);
	nand (d360, d287, d352);
	buf (d361, d299);
	buf (d362, d258);
	buf (d363, d319);
	and (d364, d276, d314);
	nand (d365, d300, d351);
	and (d366, d281, d296);
	not (d367, d158);
	nor (d368, d284, d305);
	or (d369, d307, d351);
	nand (d370, d272, d351);
	nand (d371, d286, d345);
	xor (d372, d304, d345);
	not (d373, d46);
	buf (d374, d88);
	nand (d375, d277, d306);
	not (d376, d6);
	nor (d377, d285, d327);
	buf (d378, d194);
	not (d379, d230);
	buf (d380, d308);
	nand (d381, d286, d293);
	nand (d382, d333, d347);
	nand (d383, d292, d304);
	nor (d384, d269, d302);
	nor (d385, d272, d325);
	or (d386, d331, d352);
	xor (d387, d285, d323);
	xnor (d388, d269, d320);
	xnor (d389, d310, d320);
	nand (d390, d266, d346);
	nor (d391, d301, d323);
	xnor (d392, d304, d315);
	not (d393, d282);
	and (d394, d307, d352);
	nand (d395, d327, d348);
	buf (d396, d170);
	buf (d397, d251);
	nand (d398, d300, d316);
	or (d399, d290, d299);
	and (d400, d267, d333);
	not (d401, d305);
	xor (d402, d283, d303);
	and (d403, d308, d324);
	and (d404, d333, d347);
	buf (d405, d332);
	not (d406, d303);
	nor (d407, d334, d347);
	not (d408, d299);
	buf (d409, d219);
	xor (d410, d319, d334);
	not (d411, d216);
	xor (d412, d290, d300);
	buf (d413, d161);
	not (d414, d130);
	xnor (d415, d305, d314);
	xnor (d416, d310, d334);
	nand (d417, d291, d304);
	and (d418, d286, d292);
	not (d419, d341);
	assign f1 = d381;
	assign f2 = d395;
	assign f3 = d385;
	assign f4 = d394;
endmodule
