module CCGRCG4( x0, x1, f1, f2, f3 );

	input x0, x1;
	output f1, f2, f3;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293;

	xor (d1, x1);
	not (d2, x0);
	nand (d3, x0);
	buf (d4, x1);
	nor (d5, x1);
	xor (d6, x0);
	nand (d7, x0, x1);
	buf (d8, x0);
	nand (d9, x0, x1);
	or (d10, x0, x1);
	nand (d11, x1);
	nor (d12, x0);
	or (d13, x1);
	nor (d14, x0, x1);
	xor (d15, x0, x1);
	or (d16, x0);
	or (d17, x0, x1);
	xnor (d18, x1);
	xor (d19, x0, x1);
	and (d20, x0);
	xnor (d21, x0, x1);
	xnor (d22, x0);
	not (d23, x1);
	and (d24, x1);
	xnor (d25, x0, x1);
	or (d26, d15, d18);
	or (d27, d18, d24);
	buf (d28, d15);
	nand (d29, d7, d20);
	nand (d30, d1, d13);
	and (d31, d3, d5);
	buf (d32, d14);
	nor (d33, d1, d10);
	or (d34, d6, d13);
	not (d35, d11);
	xor (d36, d3, d9);
	or (d37, d10, d14);
	and (d38, d9, d19);
	xnor (d39, d21, d23);
	or (d40, d2, d14);
	nand (d41, d16, d21);
	or (d42, d5, d8);
	nor (d43, d11, d15);
	xor (d44, d4, d10);
	nor (d45, d22, d25);
	and (d46, d3);
	and (d47, d19, d20);
	not (d48, d4);
	nor (d49, d2, d18);
	xor (d50, d12, d23);
	xor (d51, d4);
	xnor (d52, d9, d17);
	nor (d53, d4, d5);
	not (d54, d23);
	buf (d55, d21);
	xor (d56, d1, d17);
	or (d57, d13, d19);
	xnor (d58, d6, d15);
	nor (d59, d7, d11);
	nand (d60, d6, d25);
	nand (d61, d21, d23);
	xor (d62, d8, d22);
	buf (d63, d19);
	or (d64, d3, d10);
	not (d65, d1);
	not (d66, d9);
	xor (d67, d4, d16);
	and (d68, d10, d19);
	xor (d69, d7, d25);
	buf (d70, d13);
	or (d71, d3, d4);
	xor (d72, d5, d15);
	or (d73, d12, d22);
	xnor (d74, d3, d22);
	or (d75, d8, d17);
	not (d76, d25);
	or (d77, d14, d20);
	nor (d78, d22, d23);
	xnor (d79, d11, d22);
	xor (d80, d5, d8);
	xnor (d81, d16, d20);
	buf (d82, d7);
	buf (d83, d4);
	xnor (d84, d9, d14);
	xor (d85, d9, d11);
	and (d86, d11, d12);
	xnor (d87, d19);
	xor (d88, d16, d22);
	buf (d89, d11);
	nor (d90, d2, d17);
	buf (d91, d5);
	buf (d92, d22);
	not (d93, d16);
	or (d94, d7, d13);
	xnor (d95, d17, d18);
	nand (d96, d10, d12);
	xnor (d97, d14, d15);
	and (d98, d2, d8);
	xor (d99, d3, d24);
	buf (d100, d25);
	and (d101, d5, d14);
	not (d102, d19);
	and (d103, d4, d5);
	xnor (d104, d4, d6);
	nand (d105, d3, d13);
	or (d106, d2, d10);
	nor (d107, d2, d15);
	or (d108, d2, d9);
	not (d109, d5);
	nor (d110, d31, d37);
	or (d111, d64, d77);
	and (d112, d82, d100);
	not (d113, d33);
	or (d114, d56);
	or (d115, d82, d88);
	not (d116, d102);
	xnor (d117, d87, d96);
	and (d118, d64, d69);
	xnor (d119, d39, d105);
	or (d120, d63, d82);
	not (d121, d43);
	xor (d122, d28, d88);
	not (d123, d82);
	nor (d124, d26, d34);
	and (d125, d68, d89);
	xor (d126, d91, d95);
	and (d127, d86, d102);
	xnor (d128, d33, d49);
	xnor (d129, d39, d71);
	buf (d130, d104);
	not (d131, d78);
	buf (d132, d54);
	or (d133, d64, d71);
	xnor (d134, d53, d105);
	xnor (d135, d92, d109);
	and (d136, d53, d90);
	buf (d137, d105);
	or (d138, d42, d76);
	nand (d139, d38, d45);
	buf (d140, d50);
	xnor (d141, d36, d78);
	buf (d142, d3);
	or (d143, d42, d46);
	or (d144, d41, d44);
	and (d145, d38, d55);
	not (d146, d8);
	xor (d147, d28, d107);
	xnor (d148, d40, d78);
	not (d149, d51);
	or (d150, d83, d107);
	and (d151, d92, d94);
	nor (d152, d83, d109);
	or (d153, d54, d89);
	not (d154, d98);
	and (d155, d56, d102);
	xor (d156, d43, d100);
	not (d157, d39);
	or (d158, d29, d32);
	or (d159, d75, d91);
	nor (d160, d38, d73);
	and (d161, d149, d150);
	nand (d162, d132, d155);
	xor (d163, d135, d145);
	and (d164, d161, d162);
	not (d165, d68);
	xor (d166, d161, d162);
	nand (d167, d161, d162);
	nor (d168, d161, d162);
	xor (d169, d162, d163);
	nor (d170, d162, d163);
	xor (d171, d162);
	xnor (d172, d162, d163);
	nand (d173, d161, d162);
	nand (d174, d161, d163);
	or (d175, d163);
	not (d176, d65);
	xor (d177, d161, d162);
	and (d178, d161, d163);
	nor (d179, d161, d162);
	and (d180, d162, d163);
	nor (d181, d163);
	nand (d182, d161, d163);
	or (d183, d161, d162);
	xnor (d184, d161, d163);
	xnor (d185, d161);
	nor (d186, d161);
	and (d187, d163);
	not (d188, d140);
	or (d189, d162);
	buf (d190, d81);
	xnor (d191, d161, d163);
	not (d192, d12);
	buf (d193, d76);
	or (d194, d161);
	or (d195, d162, d163);
	buf (d196, d139);
	not (d197, d13);
	nor (d198, d162, d163);
	not (d199, d66);
	buf (d200, d107);
	or (d201, d161, d162);
	nand (d202, d162, d163);
	xnor (d203, d163);
	not (d204, d80);
	and (d205, d161);
	buf (d206, d41);
	buf (d207, d101);
	not (d208, d163);
	buf (d209, d118);
	xor (d210, d161);
	nand (d211, d168, d185);
	nor (d212, d208, d209);
	and (d213, d184, d194);
	nor (d214, d183, d198);
	xnor (d215, d169, d208);
	xnor (d216, d180, d192);
	nand (d217, d183, d191);
	or (d218, d166, d193);
	nor (d219, d168, d205);
	and (d220, d186, d209);
	xor (d221, d188, d196);
	not (d222, d200);
	nor (d223, d194, d198);
	not (d224, d113);
	buf (d225, d189);
	nand (d226, d181, d210);
	nor (d227, d170, d171);
	xnor (d228, d192, d198);
	nor (d229, d190, d209);
	and (d230, d186, d194);
	or (d231, d190, d192);
	or (d232, d198, d203);
	nand (d233, d178, d206);
	or (d234, d175, d193);
	buf (d235, d95);
	buf (d236, d77);
	nand (d237, d181, d183);
	not (d238, d207);
	nor (d239, d200, d207);
	nand (d240, d171, d206);
	nor (d241, d195, d199);
	nor (d242, d179, d197);
	xnor (d243, d164, d184);
	nand (d244, d179, d208);
	xnor (d245, d193, d194);
	nor (d246, d195, d198);
	and (d247, d174, d207);
	buf (d248, d48);
	buf (d249, d8);
	or (d250, d206, d210);
	nand (d251, d173, d177);
	nor (d252, d198, d200);
	nand (d253, d185, d205);
	and (d254, d167, d210);
	buf (d255, d59);
	and (d256, d166, d206);
	buf (d257, d112);
	nand (d258, d184, d187);
	or (d259, d183, d204);
	xnor (d260, d191, d210);
	not (d261, d151);
	or (d262, d190, d205);
	not (d263, d56);
	and (d264, d173);
	not (d265, d27);
	buf (d266, d69);
	nand (d267, d195, d205);
	xor (d268, d172, d181);
	not (d269, d179);
	xnor (d270, d179, d187);
	not (d271, d138);
	nand (d272, d212, d246);
	nor (d273, d211, d237);
	or (d274, d228, d234);
	buf (d275, d85);
	nand (d276, d230, d234);
	xor (d277, d236, d257);
	xor (d278, d225, d246);
	and (d279, d223, d270);
	or (d280, d215, d252);
	and (d281, d227, d256);
	or (d282, d263, d266);
	xnor (d283, d252, d256);
	nor (d284, d265, d270);
	nand (d285, d219, d261);
	and (d286, d225, d233);
	xor (d287, d213, d252);
	nand (d288, d215, d266);
	or (d289, d248, d267);
	xor (d290, d250, d268);
	nand (d291, d227, d233);
	xor (d292, d228, d246);
	xnor (d293, d228, d253);
	assign f1 = d281;
	assign f2 = d283;
	assign f3 = d290;
endmodule
