module CCGRCG12( x0, x1, f1, f2, f3, f4, f5, f6, f7 );

	input x0, x1;
	output f1, f2, f3, f4, f5, f6, f7;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304;

	nand (d1, x0, x1);
	not (d2, x0);
	or (d3, x1);
	buf (d4, x1);
	nand (d5, x1);
	xnor (d6, x0);
	buf (d7, x0);
	xor (d8, x0, x1);
	xor (d9, x1);
	xor (d10, x0);
	and (d11, x1);
	xor (d12, x0, x1);
	or (d13, d3, d5);
	xor (d14, d1, d5);
	xor (d15, d5, d7);
	not (d16, d9);
	xor (d17, d10, d12);
	nor (d18, d3, d7);
	buf (d19, d6);
	buf (d20, d12);
	xnor (d21, d8, d11);
	xor (d22, d8, d12);
	xor (d23, d7, d10);
	xnor (d24, d3, d7);
	or (d25, d1, d3);
	or (d26, d2, d6);
	not (d27, d7);
	nor (d28, d3, d10);
	buf (d29, d8);
	nand (d30, d3, d7);
	nor (d31, d1, d10);
	buf (d32, d2);
	or (d33, d3, d9);
	xnor (d34, d30);
	and (d35, d18, d32);
	xor (d36, d16, d33);
	buf (d37, d23);
	or (d38, d19, d25);
	and (d39, d21, d33);
	and (d40, d27, d29);
	and (d41, d22, d31);
	and (d42, d15, d17);
	and (d43, d19, d28);
	nand (d44, d20, d22);
	xnor (d45, d25, d29);
	and (d46, d17, d24);
	xor (d47, d16, d17);
	or (d48, d13, d15);
	nand (d49, d37, d43);
	xnor (d50, d35, d39);
	nor (d51, d41, d43);
	nor (d52, d47, d48);
	nand (d53, d50, d51);
	nor (d54, d49, d52);
	xor (d55, d51, d52);
	xor (d56, d51);
	xor (d57, d52);
	xnor (d58, d49);
	xnor (d59, d49, d50);
	and (d60, d50, d51);
	xnor (d61, d51);
	xor (d62, d50, d51);
	xnor (d63, d49, d52);
	buf (d64, d4);
	or (d65, d49, d52);
	and (d66, d49, d50);
	nand (d67, d49, d50);
	nor (d68, d51, d52);
	buf (d69, d30);
	nor (d70, d49, d51);
	not (d71, d23);
	or (d72, d50, d51);
	nand (d73, d51);
	nand (d74, d49, d50);
	and (d75, d49, d50);
	buf (d76, d18);
	xnor (d77, d50, d52);
	nor (d78, d49);
	xor (d79, d50);
	or (d80, d52);
	buf (d81, d51);
	and (d82, d49, d52);
	not (d83, d42);
	not (d84, d28);
	xor (d85, d50, d52);
	and (d86, d50, d51);
	and (d87, d52);
	and (d88, d50, d52);
	xnor (d89, d51, d52);
	xor (d90, d49, d51);
	xor (d91, d50, d52);
	not (d92, d2);
	buf (d93, d47);
	or (d94, d50, d51);
	nand (d95, d49, d51);
	xnor (d96, d49, d50);
	and (d97, d51, d52);
	nor (d98, d51, d52);
	not (d99, d13);
	xnor (d100, d49, d52);
	not (d101, d46);
	not (d102, d24);
	not (d103, d10);
	not (d104, d14);
	or (d105, d51);
	not (d106, x1);
	xnor (d107, d49, d51);
	nand (d108, d50, d52);
	nor (d109, d76, d78);
	nor (d110, d62, d63);
	nor (d111, d60, d79);
	and (d112, d76, d97);
	xor (d113, d69, d97);
	nor (d114, d89, d94);
	nand (d115, d73, d106);
	xor (d116, d70, d92);
	xnor (d117, d58, d79);
	nand (d118, d67, d72);
	nor (d119, d90, d92);
	buf (d120, d98);
	not (d121, d86);
	xnor (d122, d76, d87);
	nor (d123, d70, d78);
	xnor (d124, d82, d90);
	xor (d125, d65, d82);
	xnor (d126, d59, d83);
	nor (d127, d61, d99);
	xnor (d128, d70, d101);
	and (d129, d65, d72);
	or (d130, d86, d93);
	and (d131, d73, d80);
	xor (d132, d74, d90);
	buf (d133, d53);
	nand (d134, d78, d106);
	xor (d135, d80, d84);
	buf (d136, d20);
	buf (d137, d24);
	xor (d138, d57, d78);
	not (d139, d73);
	or (d140, d56, d107);
	or (d141, d76, d92);
	xor (d142, d73, d105);
	xor (d143, d53, d107);
	nor (d144, d80, d103);
	not (d145, d33);
	xnor (d146, d60, d90);
	xor (d147, d73, d86);
	or (d148, d69, d96);
	and (d149, d63, d89);
	not (d150, d80);
	and (d151, d69, d101);
	xnor (d152, d82, d95);
	or (d153, d60, d106);
	buf (d154, d77);
	nor (d155, d55, d58);
	and (d156, d67, d107);
	nand (d157, d74, d81);
	or (d158, d94, d99);
	or (d159, d72, d78);
	xnor (d160, d76, d77);
	xor (d161, d79, d91);
	nand (d162, d56, d107);
	xnor (d163, d54, d81);
	buf (d164, d57);
	and (d165, d79, d107);
	nand (d166, d93, d106);
	xor (d167, d71, d75);
	xnor (d168, d83, d96);
	nor (d169, d86, d97);
	buf (d170, d89);
	and (d171, d76, d94);
	xor (d172, d87, d102);
	xnor (d173, d79, d87);
	nor (d174, d58, d74);
	and (d175, d60, d81);
	and (d176, d55, d97);
	not (d177, d39);
	nand (d178, d81, d84);
	nand (d179, d57, d92);
	buf (d180, d76);
	xnor (d181, d67, d75);
	not (d182, d90);
	xor (d183, d84, d107);
	buf (d184, d31);
	nand (d185, d58, d74);
	xor (d186, d68, d80);
	or (d187, d54, d95);
	or (d188, d80, d87);
	and (d189, d81, d97);
	nor (d190, d92, d101);
	xor (d191, d72, d98);
	nand (d192, d109, d188);
	xnor (d193, d137, d190);
	xnor (d194, d123, d138);
	nor (d195, d113, d130);
	xnor (d196, d142, d160);
	or (d197, d161, d188);
	xor (d198, d140, d179);
	or (d199, d134, d155);
	nor (d200, d153, d156);
	nand (d201, d146, d157);
	and (d202, d141, d168);
	not (d203, d6);
	xor (d204, d126);
	nor (d205, d125, d160);
	and (d206, d156, d163);
	nor (d207, d123, d130);
	or (d208, d109, d174);
	buf (d209, d37);
	nand (d210, d128, d131);
	nand (d211, d132, d137);
	or (d212, d171, d183);
	or (d213, d146, d190);
	and (d214, d132, d177);
	nor (d215, d135, d168);
	xnor (d216, d111, d170);
	xor (d217, d163, d170);
	nand (d218, d141, d180);
	nand (d219, d147, d183);
	nand (d220, d134, d136);
	and (d221, d125, d161);
	or (d222, d146, d170);
	and (d223, d124, d149);
	nand (d224, d127, d148);
	nor (d225, d123, d187);
	or (d226, d145, d152);
	nand (d227, d146, d187);
	not (d228, d1);
	xor (d229, d162, d182);
	nand (d230, d139, d151);
	xnor (d231, d132, d150);
	buf (d232, d32);
	nand (d233, d141, d152);
	not (d234, d38);
	xnor (d235, d125, d131);
	or (d236, d151, d158);
	and (d237, d143, d162);
	or (d238, d119, d166);
	xor (d239, d121, d161);
	not (d240, d96);
	nand (d241, d148, d158);
	or (d242, d193, d233);
	and (d243, d209, d241);
	and (d244, d213, d236);
	and (d245, d201, d236);
	nand (d246, d195, d201);
	nor (d247, d212, d222);
	xnor (d248, d208, d209);
	xnor (d249, d231, d240);
	and (d250, d213, d223);
	buf (d251, d187);
	buf (d252, d197);
	nor (d253, d223, d235);
	nor (d254, d204, d240);
	or (d255, d208, d214);
	not (d256, d117);
	xor (d257, d201, d215);
	nor (d258, d219, d240);
	xor (d259, d206, d212);
	xnor (d260, d193, d225);
	or (d261, d238, d241);
	xor (d262, d222, d235);
	nor (d263, d206, d233);
	nand (d264, d207, d221);
	buf (d265, d188);
	nand (d266, d207, d210);
	or (d267, d195, d204);
	nor (d268, d207, d234);
	buf (d269, d68);
	and (d270, d237, d240);
	xor (d271, d195, d224);
	nor (d272, d194, d201);
	buf (d273, d148);
	nor (d274, d202, d219);
	or (d275, d196, d241);
	not (d276, d78);
	nand (d277, d230, d236);
	buf (d278, d15);
	or (d279, d205, d227);
	xnor (d280, d208, d225);
	or (d281, d201, d218);
	and (d282, d207, d241);
	nor (d283, d233, d241);
	or (d284, d211, d228);
	not (d285, d191);
	or (d286, d206, d241);
	and (d287, d221, d230);
	buf (d288, d135);
	nand (d289, d199, d222);
	and (d290, d201, d225);
	xnor (d291, d208, d214);
	nor (d292, d204, d229);
	nand (d293, d218, d241);
	not (d294, d189);
	nor (d295, d200, d234);
	and (d296, d216, d224);
	or (d297, d206, d216);
	and (d298, d201, d228);
	buf (d299, d181);
	buf (d300, d232);
	buf (d301, d227);
	nor (d302, d193, d208);
	buf (d303, d72);
	xor (d304, d205, d211);
	assign f1 = d272;
	assign f2 = d246;
	assign f3 = d271;
	assign f4 = d266;
	assign f5 = d274;
	assign f6 = d259;
	assign f7 = d291;
endmodule
