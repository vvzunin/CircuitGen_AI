module CCGRCG24( x0, x1, x2, f1, f2, f3 );

	input x0, x1, x2;
	output f1, f2, f3;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115;

	nand (d1, x1, x2);
	or (d2, x0);
	nor (d3, x0, x1);
	xnor (d4, x0, x1);
	xor (d5, x1);
	nor (d6, x1, x2);
	buf (d7, x1);
	and (d8, x2);
	not (d9, x2);
	buf (d10, x0);
	not (d11, x0);
	and (d12, x0);
	xor (d13, x0, x2);
	or (d14, x0, x1);
	nor (d15, x0, x2);
	or (d16, x1, x2);
	xor (d17, x0, x1);
	buf (d18, x2);
	and (d19, x1);
	or (d20, x0, x1);
	xnor (d21, d11, d20);
	nor (d22, d1, d19);
	nand (d23, d5, d14);
	nor (d24, d3, d6);
	nand (d25, d3, d6);
	or (d26, d10, d12);
	nand (d27, d8, d13);
	buf (d28, d13);
	or (d29, d2, d7);
	xor (d30, d18, d19);
	and (d31, d18);
	xor (d32, d2, d15);
	not (d33, x1);
	buf (d34, d20);
	xor (d35, d8, d19);
	nor (d36, d4, d14);
	or (d37, d1, d10);
	xor (d38, d7, d13);
	xor (d39, d16, d20);
	and (d40, d7, d11);
	xor (d41, d3, d11);
	nor (d42, d17, d19);
	or (d43, d6, d11);
	xnor (d44, d5, d16);
	and (d45, d1, d4);
	nand (d46, d3, d4);
	buf (d47, d4);
	xnor (d48, d13, d20);
	xnor (d49, d3, d15);
	buf (d50, d14);
	or (d51, d10, d19);
	nor (d52, d5, d14);
	and (d53, d13, d15);
	and (d54, d3, d6);
	xnor (d55, d12, d15);
	xnor (d56, d6, d16);
	nor (d57, d1, d9);
	nor (d58, d2, d8);
	xor (d59, d4, d20);
	xnor (d60, d4, d12);
	and (d61, d1, d13);
	xor (d62, d2, d13);
	not (d63, d18);
	xor (d64, d8, d9);
	buf (d65, d17);
	nor (d66, d4, d7);
	xor (d67, d13, d19);
	xor (d68, d2, d7);
	buf (d69, d11);
	or (d70, d5, d8);
	or (d71, d16);
	not (d72, d1);
	not (d73, d15);
	nand (d74, d1, d12);
	and (d75, d3, d14);
	or (d76, d1, d19);
	nand (d77, d6, d17);
	or (d78, d5, d16);
	or (d79, d2, d15);
	xor (d80, d1, d17);
	and (d81, d1, d8);
	xnor (d82, d3, d11);
	and (d83, d2, d10);
	not (d84, d55);
	or (d85, d52, d58);
	and (d86, d28, d33);
	xnor (d87, d45, d81);
	not (d88, d34);
	xor (d89, d66, d82);
	and (d90, d29, d81);
	xnor (d91, d32, d40);
	xnor (d92, d39, d50);
	and (d93, d40, d51);
	or (d94, d50, d77);
	nor (d95, d52, d74);
	not (d96, d16);
	xor (d97, d43, d66);
	or (d98, d70, d72);
	buf (d99, d69);
	xnor (d100, d55, d56);
	nor (d101, d28, d74);
	buf (d102, d77);
	nand (d103, d32, d81);
	and (d104, d41, d70);
	or (d105, d30, d65);
	or (d106, d60, d71);
	nor (d107, d25, d53);
	xnor (d108, d71, d76);
	xnor (d109, d22, d73);
	nor (d110, d38, d70);
	buf (d111, d29);
	xnor (d112, d57, d62);
	nor (d113, d58, d69);
	nor (d114, d60, d69);
	xor (d115, d56, d63);
	assign f1 = d85;
	assign f2 = d109;
	assign f3 = d84;
endmodule
