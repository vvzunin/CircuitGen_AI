module CCGRCG183( x0, x1, x2, x3, x4, x5, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17 );

	input x0, x1, x2, x3, x4, x5;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314, d315, d316, d317, d318, d319, d320, d321, d322, d323, d324, d325, d326, d327, d328, d329, d330, d331, d332, d333, d334, d335, d336, d337, d338, d339, d340, d341, d342, d343, d344, d345, d346, d347, d348, d349, d350, d351, d352, d353, d354, d355, d356, d357, d358, d359, d360, d361, d362, d363, d364, d365, d366, d367, d368, d369, d370, d371, d372, d373, d374, d375, d376, d377, d378, d379, d380, d381, d382, d383, d384, d385, d386, d387, d388, d389, d390, d391, d392, d393, d394, d395, d396, d397, d398, d399, d400, d401, d402, d403, d404, d405, d406, d407, d408, d409, d410, d411, d412, d413, d414, d415, d416, d417, d418, d419, d420, d421, d422, d423, d424, d425, d426, d427, d428, d429, d430, d431, d432, d433, d434, d435, d436, d437, d438, d439, d440, d441, d442, d443, d444, d445, d446, d447, d448, d449, d450, d451, d452, d453, d454, d455, d456, d457, d458, d459, d460, d461, d462, d463, d464, d465, d466, d467, d468, d469, d470, d471, d472, d473, d474, d475, d476, d477, d478, d479, d480, d481, d482, d483, d484, d485, d486, d487, d488, d489, d490, d491, d492, d493, d494, d495, d496, d497, d498, d499, d500, d501, d502, d503, d504, d505, d506, d507, d508, d509, d510, d511, d512, d513, d514, d515, d516, d517, d518, d519, d520, d521, d522, d523, d524, d525, d526, d527, d528, d529, d530, d531, d532, d533, d534, d535, d536, d537, d538, d539, d540, d541, d542, d543, d544, d545, d546, d547, d548, d549, d550, d551, d552, d553, d554, d555, d556, d557, d558, d559, d560, d561, d562, d563, d564, d565;

	xor (d1, x0, x3);
	buf (d2, x0);
	or (d3, x0, x1);
	or (d4, x0, x4);
	buf (d5, x3);
	xnor (d6, x2, x3);
	and (d7, x1, x5);
	and (d8, x0, x1);
	or (d9, x1, x2);
	buf (d10, x1);
	or (d11, x1, x4);
	not (d12, x5);
	xnor (d13, x3, x4);
	nor (d14, x1, x4);
	xor (d15, x3);
	and (d16, x2, x5);
	buf (d17, x5);
	and (d18, x0, x3);
	and (d19, x4, x5);
	and (d20, x2);
	not (d21, x4);
	xnor (d22, x2);
	xor (d23, x2, x3);
	nor (d24, x3, x5);
	xnor (d25, x3, x4);
	and (d26, x2, x4);
	or (d27, x3, x4);
	or (d28, x0, x5);
	nand (d29, x1, x4);
	and (d30, x1, x5);
	nand (d31, x0, x1);
	and (d32, x2, x3);
	and (d33, x1, x4);
	nor (d34, x0, x5);
	xor (d35, x0, x2);
	xnor (d36, x1);
	xor (d37, x3, x4);
	nand (d38, x0, x2);
	or (d39, x3, x5);
	and (d40, x0, x1);
	nor (d41, x4, x5);
	or (d42, x1, x3);
	xnor (d43, x0, x3);
	nand (d44, x0, x3);
	or (d45, x2);
	buf (d46, x2);
	xnor (d47, x0, x2);
	nand (d48, x0, x4);
	and (d49, x2, x3);
	buf (d50, x4);
	nand (d51, x1, x2);
	nand (d52, x4, x5);
	nor (d53, x0, x1);
	not (d54, x2);
	nand (d55, x1, x3);
	not (d56, x3);
	not (d57, x0);
	and (d58, x2, x4);
	or (d59, x4, x5);
	nand (d60, x2, x4);
	or (d61, x3);
	xnor (d62, x0, x2);
	nand (d63, x1, x2);
	nand (d64, x1, x3);
	xnor (d65, x1, x3);
	nor (d66, d9, d44);
	xor (d67, d22, d51);
	xnor (d68, d18, d20);
	nor (d69, d20, d38);
	or (d70, d31);
	not (d71, d23);
	nand (d72, d48, d54);
	xnor (d73, d30, d31);
	or (d74, d8, d26);
	buf (d75, d58);
	nand (d76, d8, d48);
	nor (d77, d15, d21);
	buf (d78, d40);
	xor (d79, d2, d31);
	buf (d80, d28);
	not (d81, d54);
	and (d82, d23, d42);
	and (d83, d9, d55);
	buf (d84, d19);
	nand (d85, d15, d36);
	buf (d86, d18);
	not (d87, d33);
	or (d88, d38, d49);
	nand (d89, d24, d49);
	xor (d90, d39, d42);
	xor (d91, d13, d16);
	buf (d92, d10);
	and (d93, d3, d38);
	nor (d94, d4, d38);
	buf (d95, d27);
	buf (d96, d46);
	buf (d97, d47);
	nand (d98, d27, d32);
	xnor (d99, d18, d52);
	xor (d100, d6, d40);
	buf (d101, d21);
	buf (d102, d41);
	not (d103, d59);
	buf (d104, d14);
	and (d105, d8, d35);
	xnor (d106, d17, d43);
	or (d107, d11, d32);
	or (d108, d4, d25);
	not (d109, d10);
	xor (d110, d10, d62);
	and (d111, d54, d59);
	xor (d112, d26, d33);
	nand (d113, d34, d39);
	nand (d114, d14, d15);
	xor (d115, d13, d59);
	nor (d116, d14, d33);
	or (d117, d48, d53);
	xnor (d118, d105, d110);
	xnor (d119, d80, d96);
	nor (d120, d71, d89);
	buf (d121, d51);
	not (d122, d40);
	xor (d123, d72, d93);
	and (d124, d85, d98);
	not (d125, d70);
	and (d126, d72, d99);
	not (d127, d73);
	not (d128, d19);
	and (d129, d74, d88);
	not (d130, d82);
	and (d131, d71, d105);
	or (d132, d125, d128);
	nand (d133, d120, d121);
	nand (d134, d127, d129);
	xor (d135, d119, d120);
	nand (d136, d123, d130);
	not (d137, d48);
	or (d138, d120, d126);
	nor (d139, d120);
	or (d140, d122, d131);
	not (d141, d6);
	xor (d142, d122, d127);
	and (d143, d118, d123);
	xor (d144, d121, d122);
	xnor (d145, d124, d127);
	and (d146, d126, d130);
	and (d147, d121, d129);
	xnor (d148, d121, d124);
	nor (d149, d121, d130);
	buf (d150, d73);
	xnor (d151, d120, d127);
	buf (d152, d92);
	not (d153, d95);
	xor (d154, d119, d127);
	buf (d155, d109);
	or (d156, d126, d127);
	xnor (d157, d122, d126);
	or (d158, d125, d129);
	nor (d159, d121, d130);
	nand (d160, d123, d129);
	xnor (d161, d120, d124);
	buf (d162, d37);
	xor (d163, d120, d128);
	xor (d164, d121, d127);
	nor (d165, d120, d128);
	xor (d166, d122, d126);
	not (d167, d74);
	not (d168, d37);
	or (d169, d127, d131);
	and (d170, d119);
	and (d171, d118, d121);
	or (d172, d126, d130);
	nor (d173, d120, d126);
	xor (d174, d121, d125);
	xor (d175, d130, d131);
	buf (d176, d114);
	buf (d177, d118);
	xor (d178, d124, d126);
	xnor (d179, d125, d128);
	not (d180, d65);
	nand (d181, d118, d121);
	buf (d182, d74);
	nor (d183, d129, d130);
	xor (d184, d123, d124);
	nor (d185, d124, d131);
	not (d186, d5);
	nand (d187, d130);
	nor (d188, d124, d126);
	and (d189, d126, d128);
	and (d190, d121, d124);
	xor (d191, d129, d130);
	xnor (d192, d120, d124);
	not (d193, d128);
	not (d194, d69);
	and (d195, d129, d130);
	or (d196, d134, d182);
	nand (d197, d154, d172);
	or (d198, d154, d191);
	or (d199, d164, d167);
	nand (d200, d163, d165);
	nand (d201, d156, d166);
	or (d202, d137, d172);
	nor (d203, d152, d164);
	nor (d204, d147, d167);
	buf (d205, d6);
	nor (d206, d162, d181);
	xor (d207, d134, d135);
	xor (d208, d143, d173);
	xor (d209, d141, d156);
	and (d210, d136, d161);
	not (d211, d28);
	or (d212, d146, d163);
	nor (d213, d134, d190);
	nor (d214, d173, d186);
	xnor (d215, d156, d191);
	and (d216, d163, d181);
	and (d217, d186, d195);
	and (d218, d155, d183);
	or (d219, d157, d187);
	nand (d220, d154, d164);
	xnor (d221, d148, d169);
	and (d222, d148, d192);
	nand (d223, d133, d151);
	nand (d224, d142, d157);
	nand (d225, d179, d193);
	nand (d226, d154, d176);
	buf (d227, d175);
	and (d228, d184);
	xor (d229, d133, d185);
	xor (d230, d153, d172);
	and (d231, d152, d182);
	xor (d232, d146, d164);
	buf (d233, d123);
	xor (d234, d177, d182);
	nand (d235, d147, d167);
	nand (d236, d155, d164);
	nor (d237, d133, d170);
	or (d238, d168, d180);
	not (d239, d31);
	or (d240, d153, d165);
	and (d241, d229, d232);
	or (d242, d211, d232);
	xor (d243, d199, d208);
	buf (d244, d185);
	and (d245, d210, d213);
	not (d246, d189);
	and (d247, d211, d232);
	not (d248, d196);
	xor (d249, d214, d224);
	nor (d250, d206, d229);
	or (d251, d215, d217);
	and (d252, d196, d210);
	xnor (d253, d201, d215);
	and (d254, d234, d235);
	not (d255, d237);
	xnor (d256, d198, d200);
	xor (d257, d196, d204);
	nor (d258, d233, d234);
	xor (d259, d227, d230);
	nand (d260, d220, d225);
	and (d261, d196, d230);
	xor (d262, d224, d239);
	nor (d263, d212, d237);
	and (d264, d211, d217);
	xor (d265, d198, d222);
	xor (d266, d200, d227);
	not (d267, d199);
	xor (d268, d230, d232);
	and (d269, d214, d219);
	or (d270, d214, d237);
	not (d271, d149);
	buf (d272, d178);
	not (d273, d143);
	not (d274, d222);
	xor (d275, d206, d229);
	xnor (d276, d218, d238);
	buf (d277, d148);
	buf (d278, d235);
	xor (d279, d202, d240);
	xor (d280, d200, d238);
	not (d281, d218);
	xor (d282, d209, d224);
	and (d283, d214, d220);
	and (d284, d211, d223);
	xor (d285, d212, d230);
	or (d286, d207, d208);
	xor (d287, d234, d235);
	xnor (d288, d213, d219);
	or (d289, d209, d210);
	or (d290, d199, d213);
	nand (d291, d200, d204);
	buf (d292, d165);
	and (d293, d217, d222);
	and (d294, d220, d224);
	not (d295, d136);
	and (d296, d224, d228);
	or (d297, d213, d236);
	xnor (d298, d225, d230);
	nand (d299, d218, d229);
	and (d300, d202, d208);
	buf (d301, d197);
	or (d302, d199, d209);
	or (d303, d215, d231);
	buf (d304, d204);
	xor (d305, d207, d237);
	nand (d306, d211, d238);
	not (d307, d51);
	not (d308, d60);
	not (d309, d216);
	xor (d310, d213, d234);
	nor (d311, d197, d224);
	xor (d312, d199, d207);
	nand (d313, d226, d232);
	or (d314, d202, d230);
	nor (d315, d218, d231);
	or (d316, d225, d227);
	xnor (d317, d198, d209);
	nor (d318, d207, d226);
	and (d319, d222, d237);
	not (d320, d44);
	nand (d321, d237, d239);
	not (d322, d111);
	or (d323, d236, d240);
	or (d324, d204, d206);
	nor (d325, d207, d219);
	nor (d326, d204, d219);
	buf (d327, d201);
	nor (d328, d241, d300);
	nor (d329, d257, d314);
	and (d330, d293, d314);
	and (d331, d277, d320);
	and (d332, d286, d307);
	and (d333, d271, d326);
	and (d334, d266, d267);
	not (d335, d232);
	xnor (d336, d307, d320);
	and (d337, d253, d256);
	not (d338, d298);
	xnor (d339, d244, d276);
	nor (d340, d289, d305);
	xnor (d341, d257, d311);
	xor (d342, d258, d316);
	nand (d343, d290, d312);
	not (d344, d224);
	nor (d345, d256, d300);
	xor (d346, d266, d326);
	buf (d347, d64);
	and (d348, d307, d312);
	or (d349, d245, d260);
	xor (d350, d256, d279);
	or (d351, d249, d294);
	xnor (d352, d268, d291);
	xor (d353, d276, d317);
	and (d354, d294, d305);
	not (d355, d266);
	and (d356, d249, d306);
	xor (d357, d287, d288);
	not (d358, d190);
	nor (d359, d253, d292);
	nand (d360, d282, d296);
	not (d361, d100);
	and (d362, d267, d319);
	and (d363, d256, d267);
	or (d364, d296, d315);
	and (d365, d244, d313);
	buf (d366, d134);
	xor (d367, d249, d325);
	nand (d368, d295, d296);
	or (d369, d290, d325);
	not (d370, d286);
	or (d371, d325, d326);
	not (d372, d205);
	xor (d373, d281, d325);
	nor (d374, d256, d316);
	xnor (d375, d258, d318);
	and (d376, d250, d293);
	not (d377, d47);
	xor (d378, d266, d305);
	nand (d379, d273, d323);
	nand (d380, d258, d276);
	not (d381, d140);
	xor (d382, d283, d314);
	and (d383, d264, d317);
	xnor (d384, d243, d251);
	xnor (d385, d254, d264);
	xnor (d386, d251, d285);
	nand (d387, d268, d289);
	nor (d388, d299, d326);
	nor (d389, d277, d290);
	xor (d390, d255, d300);
	nor (d391, d241, d249);
	or (d392, d256, d269);
	not (d393, d138);
	nand (d394, d281, d309);
	buf (d395, d93);
	nand (d396, d309, d321);
	nand (d397, d246, d270);
	xnor (d398, d258, d326);
	xnor (d399, d266, d280);
	nor (d400, d288, d314);
	or (d401, d258, d296);
	not (d402, d4);
	buf (d403, d187);
	not (d404, d67);
	not (d405, d181);
	and (d406, d276, d298);
	and (d407, d270, d278);
	nand (d408, d306, d320);
	xnor (d409, d289, d304);
	not (d410, d287);
	xnor (d411, d245, d322);
	and (d412, d338, d340);
	buf (d413, d229);
	buf (d414, d203);
	and (d415, d369, d399);
	xor (d416, d350, d369);
	not (d417, d383);
	not (d418, d281);
	buf (d419, d285);
	nand (d420, d361, d379);
	xnor (d421, d345, d409);
	nor (d422, d333, d392);
	buf (d423, d341);
	or (d424, d368, d410);
	or (d425, d370, d405);
	xnor (d426, d338, d367);
	nand (d427, d369, d379);
	and (d428, d358, d359);
	nand (d429, d348, d358);
	nor (d430, d328, d363);
	nand (d431, d400, d402);
	xor (d432, d343, d374);
	nand (d433, d403, d408);
	or (d434, d360, d411);
	xnor (d435, d349, d362);
	and (d436, d345, d393);
	xnor (d437, d330, d399);
	or (d438, d356, d374);
	xor (d439, d341, d365);
	not (d440, d393);
	or (d441, d347, d353);
	buf (d442, d236);
	buf (d443, d267);
	and (d444, d330, d348);
	xnor (d445, d336, d385);
	xnor (d446, d366, d386);
	not (d447, d248);
	and (d448, d392, d400);
	nor (d449, d383, d397);
	or (d450, d328, d387);
	xnor (d451, d365, d381);
	nor (d452, d329, d399);
	or (d453, d370, d408);
	or (d454, d333, d362);
	xnor (d455, d360, d363);
	xnor (d456, d338, d348);
	xor (d457, d375, d404);
	nand (d458, d345, d379);
	not (d459, d244);
	nor (d460, d340, d384);
	and (d461, d359, d393);
	nor (d462, d360, d380);
	nor (d463, d345, d352);
	or (d464, d393, d395);
	xnor (d465, d363, d373);
	xor (d466, d338, d364);
	or (d467, d339, d399);
	xor (d468, d338, d407);
	xnor (d469, d357, d396);
	and (d470, d356, d406);
	xor (d471, d330, d381);
	and (d472, d352, d370);
	and (d473, d335, d382);
	nor (d474, d353, d400);
	or (d475, d384, d389);
	and (d476, d380, d408);
	and (d477, d371, d406);
	and (d478, d349, d406);
	not (d479, d358);
	xor (d480, d349, d371);
	nand (d481, d333, d368);
	nor (d482, d358, d360);
	buf (d483, d306);
	nor (d484, d358, d375);
	and (d485, d371, d407);
	xnor (d486, d368, d377);
	not (d487, d132);
	xor (d488, d347, d385);
	buf (d489, d55);
	buf (d490, d206);
	and (d491, d336, d385);
	xnor (d492, d403, d410);
	nand (d493, d378, d393);
	nand (d494, d357, d389);
	nor (d495, d396, d400);
	not (d496, d274);
	buf (d497, d339);
	xnor (d498, d455, d459);
	or (d499, d425, d431);
	nand (d500, d465, d490);
	nor (d501, d463, d466);
	and (d502, d439, d472);
	buf (d503, d370);
	buf (d504, d436);
	or (d505, d423, d453);
	or (d506, d433, d480);
	nand (d507, d414, d497);
	not (d508, d352);
	xnor (d509, d450, d468);
	xor (d510, d432, d468);
	or (d511, d440, d454);
	xor (d512, d414, d456);
	xnor (d513, d442, d456);
	not (d514, d146);
	and (d515, d418, d485);
	and (d516, d412, d444);
	xnor (d517, d426, d439);
	buf (d518, d288);
	buf (d519, d176);
	nand (d520, d457, d489);
	or (d521, d451, d468);
	xor (d522, d442, d495);
	xor (d523, d428, d441);
	nor (d524, d418, d487);
	not (d525, d46);
	nand (d526, d452, d493);
	xnor (d527, d454, d479);
	xnor (d528, d460, d483);
	xor (d529, d429, d454);
	xnor (d530, d458, d463);
	nand (d531, d458, d469);
	and (d532, d434, d475);
	xnor (d533, d441, d448);
	buf (d534, d424);
	and (d535, d470, d490);
	xor (d536, d444, d485);
	or (d537, d420, d439);
	or (d538, d448, d468);
	xnor (d539, d415, d439);
	nand (d540, d414, d496);
	and (d541, d464, d488);
	nor (d542, d422, d455);
	and (d543, d447, d459);
	buf (d544, d481);
	xor (d545, d432, d478);
	xnor (d546, d449, d494);
	buf (d547, d290);
	or (d548, d443, d482);
	buf (d549, d283);
	xor (d550, d484, d485);
	or (d551, d461, d492);
	nand (d552, d449, d470);
	nor (d553, d425, d488);
	not (d554, d56);
	xnor (d555, d477, d489);
	xor (d556, d447, d449);
	nor (d557, d474, d484);
	xor (d558, d491, d492);
	xnor (d559, d442, d455);
	and (d560, d440, d441);
	nand (d561, d421, d480);
	nand (d562, d420, d440);
	and (d563, d452, d456);
	not (d564, d229);
	or (d565, d437, d438);
	assign f1 = d559;
	assign f2 = d553;
	assign f3 = d502;
	assign f4 = d507;
	assign f5 = d526;
	assign f6 = d565;
	assign f7 = d533;
	assign f8 = d506;
	assign f9 = d500;
	assign f10 = d545;
	assign f11 = d536;
	assign f12 = d556;
	assign f13 = d544;
	assign f14 = d536;
	assign f15 = d502;
	assign f16 = d513;
	assign f17 = d510;
endmodule
