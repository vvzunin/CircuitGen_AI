module CCGRCG136( x0, x1, x2, x3, x4, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13 );

	input x0, x1, x2, x3, x4;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138;

	xnor (d1, x3, x4);
	or (d2, x0, x1);
	xor (d3, x0, x1);
	nor (d4, x0, x2);
	buf (d5, x4);
	not (d6, x1);
	not (d7, x2);
	xnor (d8, x1, x4);
	nand (d9, x1, x3);
	nor (d10, x0, x1);
	xor (d11, x2, x4);
	buf (d12, x3);
	not (d13, x0);
	not (d14, x4);
	xnor (d15, x0, x1);
	nand (d16, x4);
	xnor (d17, x1, x2);
	nand (d18, x0, x1);
	xor (d19, x0);
	and (d20, x1, x4);
	nand (d21, x1);
	xor (d22, x1, x3);
	xor (d23, x1);
	xor (d24, x3, x4);
	xor (d25, x2, x4);
	nor (d26, x1, x4);
	and (d27, x2);
	or (d28, x0);
	xnor (d29, x0, x2);
	and (d30, x0);
	nand (d31, x2, x4);
	xnor (d32, x0);
	nand (d33, x0, x2);
	not (d34, x3);
	nand (d35, x0, x1);
	nor (d36, x1, x2);
	or (d37, x0, x3);
	nand (d38, x1, x2);
	xor (d39, x0, x2);
	or (d40, x1, x4);
	xor (d41, x0, x1);
	nand (d42, x2, x3);
	buf (d43, x0);
	or (d44, x0, x3);
	and (d45, x1);
	xor (d46, x1, x4);
	xor (d47, x0, x2);
	and (d48, x2, x4);
	and (d49, x0, x4);
	nand (d50, x1, x2);
	xor (d51, x1, x3);
	or (d52, x1, x3);
	nand (d53, d19, d26);
	and (d54, d11, d16);
	or (d55, d25, d44);
	xor (d56, d28, d49);
	buf (d57, d10);
	and (d58, d27, d40);
	nor (d59, d17, d29);
	nor (d60, d12, d37);
	xor (d61, d4, d12);
	or (d62, d14, d20);
	and (d63, d23, d32);
	buf (d64, d25);
	xor (d65, d47, d52);
	xnor (d66, d26, d29);
	xnor (d67, d2, d39);
	buf (d68, d2);
	and (d69, d14, d35);
	xor (d70, d13, d27);
	nand (d71, d23, d37);
	xor (d72, d7, d25);
	and (d73, d22, d38);
	and (d74, d21, d37);
	or (d75, d35, d44);
	nand (d76, d12);
	xnor (d77, d33, d47);
	buf (d78, d13);
	nor (d79, d11, d50);
	or (d80, d1, d44);
	and (d81, d19, d39);
	nor (d82, d17, d44);
	and (d83, d16, d18);
	nor (d84, d34, d46);
	nand (d85, d5, d20);
	xor (d86, d10, d22);
	buf (d87, d18);
	nor (d88, d7, d12);
	buf (d89, x2);
	not (d90, d40);
	and (d91, d4, d27);
	or (d92, d2, d23);
	and (d93, d30, d35);
	not (d94, d38);
	and (d95, d10, d12);
	not (d96, d43);
	nand (d97, d19, d34);
	or (d98, d10, d37);
	or (d99, d19, d46);
	buf (d100, d42);
	xor (d101, d3, d45);
	nor (d102, d40, d51);
	xor (d103, d20, d48);
	not (d104, d4);
	and (d105, d25, d28);
	xnor (d106, d15, d27);
	nor (d107, d20, d41);
	and (d108, d4, d26);
	xnor (d109, d9, d18);
	xnor (d110, d26, d35);
	nand (d111, d12, d44);
	xnor (d112, d3, d4);
	xor (d113, d6, d14);
	not (d114, d3);
	xor (d115, d26, d44);
	and (d116, d39);
	and (d117, d3, d46);
	buf (d118, d41);
	not (d119, d48);
	not (d120, d17);
	or (d121, d45, d52);
	nor (d122, d18, d48);
	or (d123, d9, d49);
	nor (d124, d7, d42);
	and (d125, d5, d40);
	nand (d126, d23, d24);
	nor (d127, d9, d40);
	xor (d128, d21, d25);
	not (d129, d24);
	not (d130, d1);
	xor (d131, d42);
	xnor (d132, d42, d47);
	nor (d133, d18, d32);
	not (d134, d39);
	xnor (d135, d35, d42);
	buf (d136, d48);
	or (d137, d23, d33);
	nor (d138, d20, d29);
	assign f1 = d75;
	assign f2 = d61;
	assign f3 = d64;
	assign f4 = d137;
	assign f5 = d90;
	assign f6 = d132;
	assign f7 = d53;
	assign f8 = d131;
	assign f9 = d61;
	assign f10 = d112;
	assign f11 = d67;
	assign f12 = d135;
	assign f13 = d106;
endmodule
