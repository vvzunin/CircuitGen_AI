module CCGRCG85( x0, x1, x2, x3, f1, f2, f3, f4, f5, f6 );

	input x0, x1, x2, x3;
	output f1, f2, f3, f4, f5, f6;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148;

	or (d1, x2);
	or (d2, x0, x2);
	and (d3, x2, x3);
	and (d4, x2, x3);
	xnor (d5, x1, x2);
	xnor (d6, x0, x2);
	nand (d7, x1, x2);
	or (d8, x2, x3);
	nor (d9, x2, x3);
	nor (d10, x0, x3);
	buf (d11, x0);
	nor (d12, x1, x2);
	nor (d13, x1);
	xnor (d14, x1);
	xnor (d15, x0, x2);
	nand (d16, x0, x1);
	nor (d17, x0);
	xor (d18, x0, x3);
	not (d19, x2);
	nand (d20, x0, x1);
	or (d21, x1, x3);
	xor (d22, x0, x2);
	xor (d23, x1, x3);
	xnor (d24, x1, x3);
	and (d25, x0, x3);
	xnor (d26, d4, d15);
	xnor (d27, d12, d21);
	or (d28, d3, d14);
	and (d29, d3, d11);
	buf (d30, d17);
	xnor (d31, d11, d23);
	nand (d32, d15, d17);
	and (d33, d12, d19);
	buf (d34, d15);
	or (d35, d13, d20);
	and (d36, d9, d23);
	not (d37, d5);
	not (d38, x3);
	xnor (d39, d9, d17);
	and (d40, d1, d13);
	and (d41, d6, d15);
	and (d42, d2, d14);
	buf (d43, d9);
	xor (d44, d11, d19);
	nand (d45, d2, d20);
	xor (d46, d5, d7);
	nand (d47, d13, d17);
	or (d48, d4, d23);
	not (d49, d17);
	nor (d50, d14, d15);
	nor (d51, d3, d24);
	not (d52, d13);
	nand (d53, d1, d19);
	xor (d54, d5, d12);
	xor (d55, d17, d21);
	buf (d56, d11);
	nor (d57, d30, d55);
	xor (d58, d31, d49);
	buf (d59, d47);
	nor (d60, d27, d48);
	or (d61, d29, d47);
	xor (d62, d45, d52);
	xnor (d63, d39, d46);
	or (d64, d40, d45);
	and (d65, d49, d54);
	xor (d66, d52, d56);
	or (d67, d28, d56);
	buf (d68, d10);
	nand (d69, d31, d46);
	and (d70, d53, d55);
	xnor (d71, d42, d54);
	xnor (d72, d33, d39);
	xor (d73, d37, d43);
	buf (d74, d23);
	nand (d75, d33, d47);
	nand (d76, d29, d32);
	and (d77, d38, d44);
	or (d78, d35, d39);
	xor (d79, d27, d43);
	and (d80, d30, d35);
	nor (d81, d48, d50);
	and (d82, d37, d53);
	xnor (d83, d26, d30);
	not (d84, d23);
	xor (d85, d33, d39);
	and (d86, d43, d48);
	buf (d87, d32);
	nand (d88, d30, d31);
	not (d89, d9);
	and (d90, d35, d52);
	or (d91, d35, d37);
	nand (d92, d27);
	nand (d93, d27, d54);
	buf (d94, d50);
	or (d95, d39, d43);
	xor (d96, d28, d36);
	xnor (d97, d41, d55);
	xnor (d98, d39, d52);
	nand (d99, d35, d37);
	not (d100, d39);
	buf (d101, d25);
	xor (d102, d42, d51);
	or (d103, d42, d55);
	nor (d104, d37, d50);
	nand (d105, d30, d33);
	and (d106, d28, d33);
	or (d107, d27, d36);
	buf (d108, d44);
	buf (d109, d13);
	xor (d110, d32, d35);
	xnor (d111, d33, d35);
	buf (d112, d31);
	xnor (d113, d37, d54);
	nor (d114, d31, d49);
	nor (d115, d54, d55);
	xnor (d116, d30, d44);
	nor (d117, d33, d48);
	buf (d118, d19);
	or (d119, d26, d42);
	and (d120, d29, d54);
	nor (d121, d33, d39);
	nand (d122, d27, d38);
	xnor (d123, d29, d47);
	nand (d124, d26, d31);
	not (d125, d56);
	and (d126, d45, d55);
	nor (d127, d35, d47);
	and (d128, d37, d47);
	xnor (d129, d28, d41);
	xnor (d130, d52, d54);
	xnor (d131, d37, d39);
	xnor (d132, d33, d50);
	or (d133, d30, d52);
	nor (d134, d41, d52);
	not (d135, d7);
	buf (d136, d1);
	xor (d137, d26, d45);
	xnor (d138, d40, d47);
	buf (d139, d52);
	or (d140, d46, d47);
	xnor (d141, d29, d46);
	xnor (d142, d38, d40);
	buf (d143, d49);
	xnor (d144, d33, d43);
	or (d145, d34, d53);
	nor (d146, d35, d49);
	xor (d147, d36, d52);
	xor (d148, d54, d56);
	assign f1 = d146;
	assign f2 = d92;
	assign f3 = d88;
	assign f4 = d87;
	assign f5 = d138;
	assign f6 = d104;
endmodule
