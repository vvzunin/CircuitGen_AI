module CCGRCG164( x0, x1, x2, x3, x4, x5, f1, f2, f3, f4, f5, f6, f7, f8 );

	input x0, x1, x2, x3, x4, x5;
	output f1, f2, f3, f4, f5, f6, f7, f8;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174;

	buf (d1, x0);
	nor (d2, x2, x4);
	and (d3, x0);
	and (d4, x5);
	nand (d5, x3, x5);
	xor (d6, x0, x3);
	and (d7, x2);
	xnor (d8, x2, x5);
	nand (d9, x0, x1);
	or (d10, x0, x3);
	or (d11, x0, x5);
	not (d12, x2);
	not (d13, x0);
	and (d14, x0, x5);
	not (d15, x5);
	nand (d16, x5);
	xnor (d17, x1, x2);
	buf (d18, x1);
	and (d19, x1);
	buf (d20, x2);
	xor (d21, x4);
	not (d22, x1);
	nor (d23, x2, x4);
	and (d24, x2, x3);
	nand (d25, x1, x2);
	buf (d26, x5);
	xnor (d27, x3, x5);
	not (d28, x3);
	or (d29, x3, x4);
	not (d30, x4);
	or (d31, x5);
	or (d32, x1, x3);
	xnor (d33, x0, x4);
	or (d34, x0, x1);
	or (d35, x4, x5);
	xnor (d36, x0, x5);
	xnor (d37, x1);
	nand (d38, x0);
	xnor (d39, x4);
	xnor (d40, x0);
	xnor (d41, x2);
	nor (d42, x4);
	nor (d43, x5);
	xnor (d44, x1, x4);
	xnor (d45, x1, x2);
	xnor (d46, x2, x5);
	xor (d47, x0, x5);
	and (d48, x1, x4);
	xnor (d49, x1, x5);
	nor (d50, x1, x3);
	or (d51, x1);
	xor (d52, x3, x4);
	or (d53, x0, x1);
	and (d54, x4, x5);
	or (d55, x3, x5);
	nor (d56, x2, x5);
	and (d57, x0, x4);
	or (d58, x2, x5);
	or (d59, d9);
	buf (d60, d20);
	nand (d61, d39, d42);
	buf (d62, d23);
	not (d63, d18);
	xnor (d64, d17, d47);
	xnor (d65, d5, d55);
	xnor (d66, d11, d38);
	buf (d67, d55);
	xor (d68, d12, d38);
	xor (d69, d3, d5);
	nor (d70, d48, d50);
	buf (d71, d2);
	nand (d72, d11, d36);
	xor (d73, d5, d58);
	or (d74, d17, d45);
	and (d75, d4, d17);
	nor (d76, d36, d54);
	not (d77, d24);
	or (d78, d41, d50);
	and (d79, d13, d35);
	xor (d80, d10, d22);
	and (d81, d15, d19);
	xnor (d82, d5, d40);
	nor (d83, d24, d48);
	buf (d84, d15);
	xor (d85, d27, d28);
	buf (d86, d52);
	and (d87, d15, d52);
	not (d88, d22);
	nand (d89, d23, d57);
	or (d90, d8, d23);
	nand (d91, d42, d49);
	and (d92, d10, d43);
	or (d93, d20, d31);
	or (d94, d34, d56);
	and (d95, d85, d91);
	buf (d96, d66);
	xor (d97, d79, d90);
	nand (d98, d73, d93);
	xor (d99, d80, d83);
	and (d100, d59, d85);
	xnor (d101, d64, d78);
	not (d102, d93);
	nand (d103, d82, d94);
	buf (d104, d12);
	buf (d105, d21);
	nand (d106, d80, d94);
	or (d107, d62, d89);
	nor (d108, d80, d94);
	buf (d109, d34);
	and (d110, d77, d93);
	xor (d111, d66, d94);
	nor (d112, d101, d111);
	buf (d113, d5);
	nor (d114, d95, d111);
	or (d115, d97, d98);
	nor (d116, d96, d107);
	or (d117, d104, d109);
	xnor (d118, d99, d105);
	nor (d119, d105, d107);
	not (d120, d85);
	xnor (d121, d95);
	not (d122, d94);
	nor (d123, d97, d99);
	xnor (d124, d97, d105);
	xnor (d125, d96, d100);
	buf (d126, d89);
	xnor (d127, d97, d104);
	nor (d128, d99, d110);
	and (d129, d96, d104);
	buf (d130, d9);
	xor (d131, d105, d108);
	xnor (d132, d108);
	nand (d133, d107, d108);
	xor (d134, d96, d97);
	buf (d135, d45);
	and (d136, d97);
	nor (d137, d95, d100);
	xnor (d138, d95, d106);
	or (d139, d108, d109);
	xnor (d140, d102, d104);
	buf (d141, d29);
	or (d142, d109, d110);
	not (d143, d32);
	nand (d144, d102, d105);
	or (d145, d102, d107);
	buf (d146, d35);
	nor (d147, d103, d105);
	nor (d148, d103, d105);
	nor (d149, d99, d109);
	xnor (d150, d114, d134);
	xnor (d151, d122, d144);
	and (d152, d128, d132);
	nor (d153, d124, d141);
	buf (d154, d101);
	xnor (d155, d125);
	and (d156, d125, d133);
	nand (d157, d126, d135);
	nor (d158, d128, d133);
	xnor (d159, d122, d123);
	nor (d160, d118, d142);
	xor (d161, d125, d132);
	buf (d162, d103);
	not (d163, d68);
	and (d164, d138, d145);
	xor (d165, d118, d121);
	or (d166, d123, d127);
	or (d167, d136, d138);
	xnor (d168, d121, d125);
	and (d169, d125, d149);
	xnor (d170, d116, d134);
	buf (d171, d91);
	xnor (d172, d113, d141);
	nand (d173, d145, d149);
	xnor (d174, d117, d125);
	assign f1 = d158;
	assign f2 = d151;
	assign f3 = d150;
	assign f4 = d156;
	assign f5 = d172;
	assign f6 = d160;
	assign f7 = d159;
	assign f8 = d155;
endmodule
