module CCGRCG32( x0, x1, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17, f18 );

	input x0, x1;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17, f18;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314, d315, d316, d317, d318, d319, d320, d321, d322, d323, d324, d325, d326, d327, d328, d329, d330, d331, d332, d333, d334, d335, d336, d337, d338, d339, d340, d341, d342, d343, d344, d345, d346, d347, d348, d349;

	and (d1, x0, x1);
	buf (d2, x0);
	buf (d3, x1);
	xnor (d4, x0, x1);
	nor (d5, x0);
	nand (d6, x0, x1);
	nand (d7, x1);
	not (d8, x1);
	nor (d9, x1);
	xor (d10, x0, x1);
	and (d11, x0);
	and (d12, x1);
	nand (d13, x0, x1);
	nor (d14, x0, x1);
	or (d15, x0, x1);
	or (d16, x0, x1);
	or (d17, d11, d14);
	xor (d18, d3, d15);
	and (d19, d8, d14);
	not (d20, d9);
	nand (d21, d4, d10);
	buf (d22, d6);
	not (d23, d2);
	nand (d24, d9, d16);
	xor (d25, d1, d11);
	xor (d26, d3, d5);
	or (d27, d13);
	nand (d28, d2, d16);
	nand (d29, d10, d11);
	nand (d30, d2, d11);
	xor (d31, d6, d14);
	not (d32, d14);
	not (d33, d3);
	xor (d34, d7, d9);
	xnor (d35, d9, d12);
	xnor (d36, d8, d11);
	or (d37, d6, d8);
	or (d38, d10, d16);
	buf (d39, d2);
	nor (d40, d1, d5);
	xor (d41, d1, d2);
	xor (d42, d1, d8);
	nor (d43, d4, d11);
	or (d44, d15, d16);
	buf (d45, d16);
	not (d46, d7);
	xor (d47, d16);
	nand (d48, d1, d8);
	nand (d49, d5, d16);
	nand (d50, d5, d13);
	or (d51, d4, d7);
	nor (d52, d2, d16);
	and (d53, d6, d15);
	not (d54, d8);
	xnor (d55, d1, d5);
	nand (d56, d4, d12);
	nor (d57, d2);
	or (d58, d6, d12);
	nand (d59, d2, d4);
	nand (d60, d3, d14);
	nand (d61, d1, d14);
	and (d62, d2, d10);
	and (d63, d2, d16);
	buf (d64, d15);
	xor (d65, d9, d10);
	xnor (d66, d2, d11);
	nor (d67, d20, d53);
	xnor (d68, d20, d23);
	and (d69, d37, d51);
	or (d70, d45, d62);
	and (d71, d42, d45);
	buf (d72, d65);
	nand (d73, d21, d48);
	nand (d74, d31, d42);
	not (d75, d62);
	xnor (d76, d22, d56);
	nand (d77, d19, d36);
	xor (d78, d32, d56);
	nand (d79, d36, d45);
	buf (d80, d60);
	buf (d81, d46);
	nor (d82, d24, d42);
	or (d83, d28, d36);
	not (d84, d63);
	xnor (d85, d27, d62);
	not (d86, d35);
	buf (d87, d45);
	not (d88, d26);
	nand (d89, d36, d64);
	not (d90, d59);
	and (d91, d34, d44);
	and (d92, d23, d31);
	not (d93, d64);
	or (d94, d30, d33);
	nand (d95, d53, d62);
	or (d96, d24, d45);
	buf (d97, d56);
	buf (d98, d49);
	xor (d99, d20, d54);
	buf (d100, d59);
	buf (d101, d62);
	xor (d102, d36, d48);
	or (d103, d35, d42);
	not (d104, d10);
	nor (d105, d27, d66);
	or (d106, d21, d38);
	nand (d107, d34, d61);
	xnor (d108, d22, d55);
	xnor (d109, d19, d34);
	buf (d110, d42);
	not (d111, d21);
	nor (d112, d19, d39);
	or (d113, d20, d26);
	xor (d114, d27, d49);
	or (d115, d17, d48);
	xnor (d116, d18, d48);
	buf (d117, d24);
	xnor (d118, d41, d48);
	xor (d119, d26, d40);
	xnor (d120, d29, d50);
	xor (d121, d41);
	nor (d122, d45, d60);
	and (d123, d57);
	xor (d124, d28, d32);
	nor (d125, d35, d59);
	not (d126, d11);
	or (d127, d49, d60);
	not (d128, d13);
	and (d129, d56, d60);
	not (d130, d52);
	nand (d131, d25, d28);
	not (d132, d34);
	or (d133, d21, d57);
	nor (d134, d21, d37);
	xor (d135, d56);
	or (d136, d43, d47);
	and (d137, d51, d62);
	not (d138, d65);
	not (d139, d41);
	xor (d140, d24, d45);
	xor (d141, d24, d35);
	nand (d142, d17, d26);
	not (d143, d15);
	nor (d144, d19, d43);
	nand (d145, d19, d32);
	nor (d146, d39, d58);
	xnor (d147, d32, d47);
	xnor (d148, d23, d31);
	nor (d149, d28, d40);
	and (d150, d32, d39);
	xor (d151, d28, d53);
	and (d152, d33, d55);
	xor (d153, d39, d63);
	xor (d154, d48, d63);
	not (d155, d113);
	or (d156, d90, d150);
	buf (d157, d148);
	nor (d158, d79, d138);
	not (d159, d19);
	not (d160, d4);
	not (d161, d88);
	nand (d162, d85, d96);
	not (d163, d120);
	and (d164, d109, d110);
	nor (d165, d158, d159);
	or (d166, d157, d162);
	nor (d167, d155, d161);
	or (d168, d163);
	nand (d169, d159, d162);
	not (d170, d67);
	or (d171, d161, d164);
	xor (d172, d156, d159);
	nand (d173, d155, d164);
	buf (d174, d101);
	nand (d175, d160);
	buf (d176, d85);
	buf (d177, d119);
	xnor (d178, d158);
	xor (d179, d159, d162);
	not (d180, d30);
	xor (d181, d158, d161);
	and (d182, d155, d164);
	xnor (d183, d160, d163);
	buf (d184, d29);
	nor (d185, d158, d163);
	buf (d186, d90);
	and (d187, d158, d162);
	xnor (d188, d159, d162);
	or (d189, d155, d157);
	buf (d190, d25);
	not (d191, d16);
	or (d192, d158, d160);
	xnor (d193, d155, d161);
	nor (d194, d160, d164);
	nor (d195, d160, d163);
	or (d196, d162, d163);
	xor (d197, d161, d162);
	buf (d198, d33);
	xor (d199, d158, d164);
	nand (d200, d161, d163);
	nor (d201, d158, d162);
	and (d202, d155, d156);
	nor (d203, d159, d164);
	xnor (d204, d157, d159);
	nor (d205, d155);
	not (d206, d140);
	and (d207, d155, d163);
	and (d208, d157, d164);
	or (d209, d155);
	xor (d210, d155, d164);
	xnor (d211, d160, d164);
	not (d212, d87);
	xor (d213, d160, d164);
	not (d214, d142);
	xor (d215, d155, d161);
	buf (d216, d94);
	or (d217, d158, d161);
	and (d218, d160, d164);
	nor (d219, d156);
	and (d220, d161, d163);
	nand (d221, d158, d161);
	not (d222, d163);
	nor (d223, d157, d160);
	and (d224, d159, d164);
	not (d225, d96);
	nor (d226, d157, d164);
	nand (d227, d156, d157);
	not (d228, d81);
	not (d229, d114);
	or (d230, d156, d158);
	and (d231, d155, d162);
	xnor (d232, d157, d161);
	nand (d233, d160, d162);
	buf (d234, d116);
	nor (d235, d162, d164);
	or (d236, d158, d159);
	xnor (d237, d156, d163);
	xnor (d238, d160, d163);
	buf (d239, d37);
	or (d240, d156, d157);
	and (d241, d158, d161);
	not (d242, d129);
	and (d243, d161, d162);
	and (d244, d159, d163);
	buf (d245, d67);
	nor (d246, d159, d163);
	xor (d247, d159);
	nor (d248, d156, d164);
	nand (d249, d157, d159);
	nor (d250, d158, d160);
	and (d251, d155, d158);
	and (d252, d158, d160);
	buf (d253, d72);
	or (d254, d155, d160);
	nor (d255, d157, d160);
	xnor (d256, d155, d164);
	buf (d257, d53);
	nand (d258, d167, d218);
	nor (d259, d167, d214);
	and (d260, d194, d246);
	xnor (d261, d249, d254);
	xnor (d262, d201, d246);
	nand (d263, d197, d211);
	or (d264, d174, d200);
	xor (d265, d170, d180);
	buf (d266, d144);
	xnor (d267, d166, d200);
	xnor (d268, d183, d221);
	or (d269, d234, d249);
	or (d270, d171, d246);
	buf (d271, d216);
	xnor (d272, d202, d243);
	buf (d273, d13);
	nor (d274, d242, d256);
	buf (d275, d111);
	or (d276, d225, d251);
	and (d277, d205, d254);
	nand (d278, d176, d185);
	or (d279, d214, d221);
	xor (d280, d175, d243);
	nand (d281, d225, d242);
	and (d282, d209, d234);
	or (d283, d191, d206);
	xnor (d284, d206, d242);
	nand (d285, d192, d241);
	xnor (d286, d189, d213);
	nor (d287, d221, d254);
	and (d288, d181, d250);
	nor (d289, d187, d225);
	nand (d290, d196, d198);
	xor (d291, d196, d232);
	buf (d292, d117);
	nand (d293, d165, d175);
	xor (d294, d179, d225);
	or (d295, d167, d215);
	xnor (d296, d182, d199);
	nand (d297, d194, d218);
	and (d298, d230, d236);
	nand (d299, d192, d199);
	xor (d300, d171, d188);
	nand (d301, d223, d249);
	xor (d302, d202, d243);
	xor (d303, d205, d229);
	buf (d304, d135);
	nor (d305, d259, d266);
	nor (d306, d286, d303);
	nor (d307, d273, d286);
	nand (d308, d273, d289);
	nand (d309, d260, d285);
	buf (d310, d247);
	not (d311, d228);
	or (d312, d284, d286);
	nor (d313, d278, d287);
	buf (d314, d300);
	xnor (d315, d263, d288);
	xnor (d316, d273, d297);
	not (d317, d155);
	buf (d318, d282);
	nor (d319, d281, d304);
	not (d320, x0);
	nand (d321, d257, d291);
	xor (d322, d261, d299);
	not (d323, d225);
	nand (d324, d259, d298);
	buf (d325, d193);
	or (d326, d282, d296);
	and (d327, d258, d284);
	or (d328, d264, d286);
	or (d329, d266, d291);
	not (d330, d27);
	nand (d331, d268, d272);
	nor (d332, d296, d297);
	and (d333, d275, d295);
	xor (d334, d287, d297);
	or (d335, d295, d297);
	not (d336, d289);
	not (d337, d109);
	nand (d338, d287, d291);
	nor (d339, d265, d281);
	nand (d340, d260, d289);
	nand (d341, d277, d278);
	or (d342, d280, d285);
	or (d343, d267, d304);
	or (d344, d263, d271);
	nand (d345, d257, d297);
	buf (d346, d202);
	and (d347, d302, d303);
	not (d348, d82);
	and (d349, d291, d302);
	assign f1 = d345;
	assign f2 = d346;
	assign f3 = d313;
	assign f4 = d319;
	assign f5 = d340;
	assign f6 = d347;
	assign f7 = d333;
	assign f8 = d317;
	assign f9 = d347;
	assign f10 = d316;
	assign f11 = d325;
	assign f12 = d307;
	assign f13 = d312;
	assign f14 = d319;
	assign f15 = d344;
	assign f16 = d342;
	assign f17 = d346;
	assign f18 = d340;
endmodule
