module CCGRCG12( x0, x1, f1, f2, f3, f4, f5, f6, f7, f8 );

	input x0, x1;
	output f1, f2, f3, f4, f5, f6, f7, f8;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314, d315, d316, d317, d318, d319, d320, d321, d322, d323, d324, d325, d326, d327, d328, d329, d330, d331, d332, d333, d334, d335, d336, d337, d338, d339, d340, d341, d342, d343, d344, d345, d346, d347, d348, d349, d350, d351, d352, d353, d354, d355, d356, d357, d358, d359, d360, d361, d362, d363, d364, d365, d366, d367, d368, d369, d370, d371, d372, d373, d374, d375, d376, d377, d378, d379, d380, d381, d382, d383, d384, d385, d386, d387, d388, d389, d390, d391, d392, d393, d394, d395, d396, d397, d398, d399, d400, d401, d402, d403, d404, d405, d406, d407, d408, d409, d410, d411, d412, d413, d414, d415, d416, d417, d418, d419, d420, d421, d422, d423, d424, d425, d426, d427, d428, d429, d430, d431, d432, d433, d434, d435, d436, d437, d438, d439, d440, d441, d442;

	buf (d1, x1);
	nand (d2, x1);
	xor (d3, x1);
	and (d4, x0, x1);
	buf (d5, x0);
	xor (d6, x0, x1);
	nor (d7, x0, x1);
	nand (d8, x0, x1);
	nand (d9, x0, x1);
	nor (d10, x0);
	or (d11, x0, x1);
	nor (d12, x1);
	or (d13, x0);
	nor (d14, x0, x1);
	xor (d15, x0, x1);
	not (d16, x1);
	not (d17, x0);
	or (d18, x0, x1);
	or (d19, x1);
	and (d20, x0);
	nand (d21, x0);
	xnor (d22, x0, x1);
	xor (d23, x0);
	and (d24, x0, x1);
	and (d25, x1);
	xnor (d26, x1);
	xor (d27, d17, d24);
	not (d28, d12);
	xor (d29, d5, d9);
	not (d30, d20);
	xor (d31, d7, d10);
	nand (d32, d13, d20);
	xor (d33, d13, d14);
	buf (d34, d17);
	xor (d35, d13, d17);
	buf (d36, d10);
	buf (d37, d12);
	or (d38, d21, d25);
	buf (d39, d9);
	and (d40, d1, d8);
	nand (d41, d22, d25);
	buf (d42, d19);
	buf (d43, d4);
	and (d44, d1, d3);
	xnor (d45, d25, d26);
	buf (d46, d13);
	or (d47, d4, d8);
	or (d48, d4, d15);
	and (d49, d17, d18);
	xnor (d50, d3, d20);
	nand (d51, d3, d16);
	buf (d52, d1);
	or (d53, d2, d20);
	nand (d54, d12, d16);
	xor (d55, d5, d20);
	xnor (d56, d8);
	or (d57, d7, d15);
	or (d58, d4, d14);
	nand (d59, d14, d25);
	xnor (d60, d8, d25);
	xnor (d61, d20, d24);
	buf (d62, d7);
	nor (d63, d1, d3);
	nor (d64, d15, d26);
	buf (d65, d23);
	xor (d66, d2, d21);
	or (d67, d11, d12);
	buf (d68, d11);
	xor (d69, d19, d23);
	nor (d70, d3, d22);
	not (d71, d10);
	or (d72, d7, d24);
	xor (d73, d10, d15);
	nand (d74, d17, d22);
	xor (d75, d3);
	buf (d76, d6);
	nand (d77, d4, d5);
	xnor (d78, d10, d21);
	and (d79, d2, d6);
	nand (d80, d7, d20);
	xnor (d81, d2, d9);
	nor (d82, d12, d16);
	nand (d83, d4, d23);
	nor (d84, d9);
	not (d85, d4);
	not (d86, d9);
	nand (d87, d1, d11);
	xor (d88, d11, d18);
	not (d89, d46);
	xnor (d90, d51, d75);
	buf (d91, d20);
	xor (d92, d37, d82);
	not (d93, d64);
	xor (d94, d30, d74);
	not (d95, d66);
	xor (d96, d47, d64);
	not (d97, d29);
	nor (d98, d44, d46);
	xnor (d99, d44, d84);
	nand (d100, d31);
	and (d101, d58, d87);
	xor (d102, d53, d83);
	and (d103, d45, d54);
	and (d104, d51, d88);
	nor (d105, d62, d77);
	xor (d106, d65, d82);
	and (d107, d29, d40);
	buf (d108, d41);
	not (d109, d53);
	nor (d110, d34, d66);
	and (d111, d51, d66);
	nor (d112, d31, d72);
	xnor (d113, d39, d67);
	nor (d114, d34, d65);
	nand (d115, d30, d85);
	xnor (d116, d45, d53);
	nor (d117, d43, d49);
	nor (d118, d65, d88);
	or (d119, d69, d80);
	buf (d120, d18);
	buf (d121, d26);
	xnor (d122, d31, d57);
	xnor (d123, d68, d78);
	nor (d124, d45, d63);
	not (d125, d55);
	and (d126, d66, d81);
	nand (d127, d35, d40);
	and (d128, d42, d43);
	or (d129, d36, d68);
	and (d130, d50, d68);
	and (d131, d36, d48);
	xnor (d132, d30, d46);
	not (d133, d23);
	nand (d134, d100, d116);
	xor (d135, d102, d106);
	buf (d136, d74);
	xnor (d137, d105, d116);
	xor (d138, d108, d118);
	nand (d139, d92, d106);
	or (d140, d95, d107);
	xnor (d141, d116, d119);
	or (d142, d89, d108);
	buf (d143, d111);
	buf (d144, d104);
	buf (d145, d93);
	nor (d146, d114, d127);
	xor (d147, d118, d132);
	or (d148, d95, d98);
	buf (d149, d79);
	and (d150, d129, d132);
	xnor (d151, d90, d114);
	nor (d152, d93, d112);
	buf (d153, d87);
	nand (d154, d93, d112);
	nand (d155, d93, d127);
	xnor (d156, d112, d126);
	xnor (d157, d128);
	nand (d158, d102, d129);
	xor (d159, d89, d105);
	buf (d160, d37);
	nand (d161, d93, d116);
	nor (d162, d100, d132);
	buf (d163, d36);
	nor (d164, d116, d131);
	buf (d165, d89);
	or (d166, d90, d128);
	nor (d167, d110, d129);
	nor (d168, d105, d107);
	xnor (d169, d99, d105);
	buf (d170, d84);
	xnor (d171, d99, d108);
	not (d172, d124);
	nor (d173, d106, d123);
	nand (d174, d90, d105);
	not (d175, d102);
	xnor (d176, d114);
	nor (d177, d115, d116);
	not (d178, d105);
	not (d179, d80);
	and (d180, d97, d128);
	not (d181, d15);
	nand (d182, d106, d108);
	and (d183, d110, d112);
	nand (d184, d91, d115);
	buf (d185, d28);
	nor (d186, d141, d180);
	and (d187, d156, d176);
	or (d188, d178, d181);
	xnor (d189, d147, d183);
	buf (d190, d25);
	or (d191, d161, d179);
	xnor (d192, d159, d183);
	nor (d193, d153, d165);
	or (d194, d162, d166);
	xor (d195, d135, d155);
	or (d196, d136, d170);
	buf (d197, d99);
	xor (d198, d139, d164);
	buf (d199, d137);
	and (d200, d166, d176);
	nor (d201, d148, d179);
	or (d202, d145, d181);
	not (d203, d96);
	xor (d204, d133, d160);
	and (d205, d174, d179);
	xnor (d206, d135, d151);
	and (d207, d147, d163);
	nand (d208, d145, d156);
	nand (d209, d133, d176);
	buf (d210, d62);
	nand (d211, d154, d161);
	and (d212, d134, d146);
	xor (d213, d142, d168);
	and (d214, d165, d176);
	not (d215, d177);
	nor (d216, d140, d142);
	xnor (d217, d157);
	and (d218, d141, d185);
	xor (d219, d159, d172);
	nand (d220, d159, d171);
	not (d221, d114);
	nand (d222, d139, d155);
	nand (d223, d169, d171);
	and (d224, d147, d155);
	or (d225, d163, d173);
	and (d226, d140, d163);
	nor (d227, d155, d175);
	xor (d228, d137, d179);
	nor (d229, d172, d181);
	xor (d230, d139, d174);
	nand (d231, d225, d228);
	not (d232, d37);
	nor (d233, d195, d211);
	or (d234, d215, d217);
	xnor (d235, d186, d201);
	not (d236, d132);
	xnor (d237, d192, d220);
	nor (d238, d191, d211);
	xnor (d239, d206, d214);
	nor (d240, d205, d208);
	xnor (d241, d202, d203);
	and (d242, d196, d221);
	xor (d243, d194, d219);
	xor (d244, d218, d222);
	or (d245, d192, d205);
	nand (d246, d188, d228);
	or (d247, d211, d219);
	or (d248, d198, d204);
	xor (d249, d191, d194);
	and (d250, d198, d209);
	nand (d251, d199, d219);
	nand (d252, d201, d203);
	buf (d253, d69);
	or (d254, d187, d228);
	nor (d255, d195, d217);
	xor (d256, d216, d219);
	xor (d257, d186, d228);
	nor (d258, d201, d228);
	and (d259, d201, d230);
	nor (d260, d188, d212);
	not (d261, d178);
	nor (d262, d188, d230);
	or (d263, d188, d209);
	xnor (d264, d196, d201);
	xor (d265, d197, d226);
	not (d266, d182);
	nor (d267, d191, d213);
	xor (d268, d193, d214);
	nor (d269, d210, d214);
	nand (d270, d203, d225);
	and (d271, d203);
	or (d272, d193, d194);
	xor (d273, d195, d208);
	xor (d274, d188, d193);
	and (d275, d196, d208);
	xnor (d276, d215, d229);
	nand (d277, d192, d221);
	nor (d278, d215, d219);
	or (d279, d188, d221);
	nand (d280, d210, d224);
	nor (d281, d194, d202);
	not (d282, d75);
	or (d283, d192, d195);
	or (d284, d196, d204);
	or (d285, d188, d222);
	xor (d286, d216, d220);
	and (d287, d204, d226);
	buf (d288, d130);
	and (d289, d186, d228);
	xor (d290, d210, d216);
	xnor (d291, d218, d219);
	buf (d292, d115);
	nor (d293, d223, d226);
	nand (d294, d210, d218);
	xor (d295, d189, d220);
	xnor (d296, d212, d230);
	xnor (d297, d222, d225);
	or (d298, d193, d209);
	nand (d299, d190, d227);
	not (d300, d98);
	nand (d301, d216, d227);
	xor (d302, d219, d221);
	or (d303, d199, d221);
	nand (d304, d198, d229);
	buf (d305, d34);
	xor (d306, d192, d196);
	xnor (d307, d190, d203);
	and (d308, d211, d219);
	xor (d309, d199, d218);
	xor (d310, d201, d217);
	nor (d311, d202, d207);
	and (d312, d199, d211);
	and (d313, d205, d227);
	not (d314, d45);
	buf (d315, d117);
	not (d316, d60);
	or (d317, d190, d194);
	buf (d318, d73);
	xnor (d319, d196, d213);
	not (d320, d187);
	buf (d321, d233);
	buf (d322, d275);
	or (d323, d263, d273);
	nand (d324, d231, d307);
	nand (d325, d278, d295);
	not (d326, d32);
	nor (d327, d244, d258);
	buf (d328, d116);
	nor (d329, d272, d309);
	nand (d330, d250, d275);
	or (d331, d259, d306);
	not (d332, d259);
	and (d333, d244, d254);
	nor (d334, d238, d269);
	xor (d335, d260, d269);
	xnor (d336, d242, d280);
	xnor (d337, d251, d294);
	or (d338, d284, d294);
	buf (d339, d120);
	nand (d340, d259, d263);
	or (d341, d235, d251);
	xor (d342, d306, d312);
	not (d343, d120);
	nand (d344, d245, d248);
	and (d345, d235, d302);
	xnor (d346, d259, d292);
	nand (d347, d297, d305);
	and (d348, d232, d258);
	xor (d349, d286, d320);
	nand (d350, d251, d319);
	nand (d351, d273, d303);
	not (d352, d65);
	nand (d353, d266, d267);
	xor (d354, d253, d263);
	not (d355, d223);
	not (d356, d116);
	xor (d357, d257, d261);
	xnor (d358, d251, d311);
	nor (d359, d274, d281);
	xnor (d360, d246, d302);
	and (d361, d247, d275);
	xnor (d362, d268, d280);
	nor (d363, d251, d308);
	and (d364, d237, d289);
	and (d365, d276, d309);
	nor (d366, d235, d271);
	buf (d367, d106);
	xnor (d368, d259, d274);
	and (d369, d250, d310);
	xor (d370, d282, d319);
	xnor (d371, d318);
	xor (d372, d277, d316);
	not (d373, d137);
	or (d374, d235, d314);
	xor (d375, d262, d273);
	xor (d376, d234, d295);
	buf (d377, d163);
	or (d378, d238, d241);
	buf (d379, d71);
	and (d380, d254, d301);
	xor (d381, d243, d299);
	xnor (d382, d257, d288);
	buf (d383, d131);
	xnor (d384, d276, d309);
	nor (d385, d236, d265);
	nor (d386, d267, d283);
	nor (d387, d262, d306);
	buf (d388, d77);
	xor (d389, d277);
	buf (d390, d237);
	xnor (d391, d347, d390);
	nor (d392, d348, d360);
	xor (d393, d345, d390);
	and (d394, d327, d331);
	buf (d395, d280);
	nor (d396, d349, d358);
	or (d397, d341, d352);
	nand (d398, d324, d381);
	buf (d399, d328);
	nor (d400, d340, d349);
	xor (d401, d357, d385);
	xnor (d402, d325, d372);
	or (d403, d364, d365);
	xor (d404, d348, d362);
	nor (d405, d323, d375);
	xor (d406, d324, d355);
	and (d407, d327, d359);
	xnor (d408, d368, d379);
	xor (d409, d339, d354);
	nand (d410, d333, d375);
	nand (d411, d329, d388);
	xnor (d412, d344, d355);
	or (d413, d367, d379);
	xnor (d414, d333, d373);
	nor (d415, d327, d390);
	or (d416, d325, d352);
	or (d417, d360, d384);
	xnor (d418, d326, d339);
	nand (d419, d346, d379);
	xor (d420, d344, d363);
	xnor (d421, d363, d379);
	nor (d422, d353, d376);
	buf (d423, d108);
	nand (d424, d334, d382);
	not (d425, d230);
	not (d426, d113);
	xor (d427, d343, d352);
	and (d428, d345, d360);
	and (d429, d336, d342);
	xnor (d430, d358, d362);
	and (d431, d363, d378);
	buf (d432, d154);
	buf (d433, d362);
	xor (d434, d335, d355);
	or (d435, d334, d349);
	nor (d436, d323, d356);
	and (d437, d332, d353);
	xnor (d438, d350, d371);
	buf (d439, d241);
	xnor (d440, d339, d372);
	or (d441, d340, d364);
	buf (d442, d24);
	assign f1 = d436;
	assign f2 = d423;
	assign f3 = d404;
	assign f4 = d429;
	assign f5 = d439;
	assign f6 = d391;
	assign f7 = d406;
	assign f8 = d435;
endmodule
