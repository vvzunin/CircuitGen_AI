// Benchmark "CCGRCG48" written by ABC on Tue Feb 13 20:51:37 2024

module CCGRCG48 ( 
    x0, x1, x2,
    f1, f2, f3, f4, f5, f6, f7  );
  input  x0, x1, x2;
  output f1, f2, f3, f4, f5, f6, f7;
  assign f1 = ~x0;
  assign f2 = ~x0 & ~x2;
  assign f3 = x1 & x2;
  assign f6 = ~x1;
  assign f4 = ~x0 & ~x2;
  assign f5 = ~x0;
  assign f7 = x1 & x2;
endmodule


