module CCGRCG191( x0, x1, x2, x3, x4, x5, x6, f1, f2 );

	input x0, x1, x2, x3, x4, x5, x6;
	output f1, f2;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250;

	or (d1, x0, x6);
	not (d2, x3);
	buf (d3, x4);
	nand (d4, x1, x2);
	nor (d5, x5);
	nor (d6, x6);
	nor (d7, x3, x5);
	nor (d8, x4);
	nor (d9, x1, x6);
	and (d10, x3, x5);
	xor (d11, x5, x6);
	and (d12, x0, x5);
	not (d13, x1);
	buf (d14, x0);
	buf (d15, x1);
	nand (d16, x2, x3);
	or (d17, x2, x4);
	or (d18, x0, x5);
	not (d19, x0);
	and (d20, x4);
	xnor (d21, x0, x5);
	and (d22, x1, x2);
	xor (d23, x2, x6);
	nand (d24, x3, x5);
	buf (d25, x2);
	and (d26, x1, x4);
	xnor (d27, x2, x4);
	or (d28, x2, x4);
	buf (d29, x3);
	xor (d30, x2);
	nor (d31, x1, x5);
	xnor (d32, x1, x6);
	xnor (d33, x4);
	or (d34, x0, x2);
	and (d35, x0, x6);
	xnor (d36, x6);
	or (d37, x1, x3);
	and (d38, x3, x5);
	xor (d39, x1, x3);
	not (d40, x5);
	nand (d41, x0, x5);
	or (d42, x0, x1);
	xor (d43, x0, x5);
	nor (d44, x5, x6);
	nand (d45, x6);
	nor (d46, x2, x5);
	buf (d47, x6);
	nand (d48, x0, x3);
	or (d49, x0, x5);
	buf (d50, d10);
	not (d51, d29);
	nand (d52, d36, d40);
	xor (d53, d26, d49);
	xnor (d54, d15, d33);
	buf (d55, d33);
	buf (d56, d47);
	xnor (d57, d18, d27);
	xnor (d58, d19, d27);
	nor (d59, d18, d36);
	xnor (d60, d36, d38);
	and (d61, d42, d46);
	or (d62, d10, d17);
	or (d63, d3, d38);
	buf (d64, d31);
	xnor (d65, d9, d14);
	xnor (d66, d1, d17);
	nor (d67, d1, d7);
	not (d68, d8);
	nand (d69, d12, d31);
	or (d70, d13, d44);
	not (d71, d3);
	not (d72, d25);
	xnor (d73, d5, d49);
	not (d74, d42);
	and (d75, d3, d28);
	nor (d76, d10, d31);
	and (d77, d10, d37);
	and (d78, d18, d34);
	nor (d79, d25, d46);
	buf (d80, d48);
	buf (d81, d19);
	buf (d82, d15);
	not (d83, d1);
	nand (d84, d35, d42);
	nand (d85, d30, d36);
	or (d86, d29, d48);
	xnor (d87, d37, d42);
	or (d88, d20, d31);
	buf (d89, d4);
	not (d90, d44);
	xnor (d91, d19, d38);
	or (d92, d22, d35);
	buf (d93, d11);
	xnor (d94, d4, d12);
	xor (d95, d7, d27);
	xor (d96, d12, d33);
	buf (d97, d45);
	xnor (d98, d29, d30);
	nand (d99, d6, d42);
	not (d100, d24);
	or (d101, d11, d12);
	xnor (d102, d13, d37);
	not (d103, d35);
	nor (d104, d18, d38);
	or (d105, d23, d43);
	xor (d106, d10, d47);
	not (d107, d75);
	not (d108, d41);
	or (d109, d74, d104);
	nor (d110, d57, d106);
	nand (d111, d68, d72);
	xor (d112, d66, d103);
	or (d113, d84, d101);
	nand (d114, d76, d82);
	buf (d115, d99);
	nand (d116, d53, d73);
	xor (d117, d72, d98);
	nand (d118, d53, d89);
	nand (d119, d55, d92);
	nand (d120, d86, d105);
	not (d121, d7);
	xnor (d122, d50, d68);
	and (d123, d58, d77);
	xnor (d124, d92, d97);
	xnor (d125, d87, d96);
	xor (d126, d62, d101);
	nor (d127, d52, d98);
	xnor (d128, d78, d81);
	not (d129, d53);
	buf (d130, d3);
	nand (d131, d83, d84);
	buf (d132, d106);
	xor (d133, d58, d67);
	nand (d134, d51, d73);
	nor (d135, d51, d100);
	xnor (d136, d70, d99);
	nor (d137, d85, d106);
	xor (d138, d61, d103);
	or (d139, d64, d88);
	not (d140, d9);
	xnor (d141, d59, d61);
	xor (d142, d72, d96);
	buf (d143, d74);
	buf (d144, d92);
	nor (d145, d67, d78);
	xor (d146, d75, d77);
	xor (d147, d74, d92);
	or (d148, d80, d93);
	xor (d149, d57, d59);
	not (d150, d104);
	xor (d151, d75, d105);
	buf (d152, d72);
	buf (d153, d13);
	not (d154, d98);
	and (d155, d55, d89);
	and (d156, d86, d96);
	xor (d157, d51, d70);
	nand (d158, d63, d91);
	or (d159, d67, d96);
	buf (d160, d57);
	nor (d161, d63, d98);
	xor (d162, d87, d94);
	or (d163, d71, d87);
	nor (d164, d64, d98);
	nor (d165, d73, d84);
	xnor (d166, d73, d94);
	xnor (d167, d56, d74);
	nor (d168, d59, d67);
	not (d169, x6);
	buf (d170, d97);
	nand (d171, d68, d96);
	buf (d172, d32);
	xnor (d173, d69, d88);
	not (d174, d31);
	and (d175, d77, d104);
	or (d176, d130, d150);
	or (d177, d153, d159);
	buf (d178, d77);
	not (d179, d155);
	xor (d180, d155, d175);
	xnor (d181, d140, d155);
	xor (d182, d134, d168);
	nand (d183, d117, d137);
	buf (d184, d43);
	nor (d185, d123, d160);
	not (d186, d174);
	or (d187, d128, d148);
	and (d188, d123, d150);
	or (d189, d148, d163);
	or (d190, d116, d169);
	nand (d191, d130, d162);
	xnor (d192, d108, d134);
	not (d193, d167);
	buf (d194, x5);
	nand (d195, d116, d145);
	or (d196, d156, d171);
	or (d197, d167, d171);
	or (d198, d115, d138);
	not (d199, d50);
	xor (d200, d124, d138);
	or (d201, d134, d174);
	xnor (d202, d131, d144);
	nand (d203, d128, d149);
	and (d204, d116, d159);
	and (d205, d131, d142);
	xnor (d206, d132, d175);
	and (d207, d139, d144);
	buf (d208, d113);
	and (d209, d128, d160);
	xor (d210, d151, d154);
	nor (d211, d153, d169);
	xnor (d212, d122, d138);
	xor (d213, d120, d167);
	buf (d214, d146);
	and (d215, d156, d173);
	nand (d216, d133, d145);
	and (d217, d131, d162);
	and (d218, d119, d168);
	nand (d219, d158, d165);
	xnor (d220, d139, d159);
	buf (d221, d118);
	xnor (d222, d134, d156);
	or (d223, d165, d174);
	nor (d224, d132, d168);
	and (d225, d129, d160);
	nand (d226, d111, d150);
	and (d227, d132, d171);
	nand (d228, d144, d171);
	xnor (d229, d131, d152);
	or (d230, d110, d159);
	xnor (d231, d167, d172);
	xnor (d232, d128, d135);
	not (d233, d45);
	xnor (d234, d112, d129);
	xnor (d235, d120, d140);
	nor (d236, d153, d158);
	nand (d237, d112, d138);
	or (d238, d147, d160);
	and (d239, d119, d131);
	nand (d240, d132, d161);
	not (d241, d94);
	xnor (d242, d142, d170);
	xnor (d243, d108, d118);
	buf (d244, d88);
	xnor (d245, d130, d162);
	buf (d246, d39);
	nand (d247, d114, d147);
	nand (d248, d125, d164);
	nor (d249, d136, d149);
	or (d250, d124, d127);
	assign f1 = d250;
	assign f2 = d237;
endmodule
