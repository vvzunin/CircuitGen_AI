module CCGRCG8( x0, x1, f1, f2, f3, f4, f5 );

	input x0, x1;
	output f1, f2, f3, f4, f5;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143;

	or (d1, x1);
	nand (d2, x0, x1);
	buf (d3, x0);
	nand (d4, x0);
	or (d5, d1, d3);
	nor (d6, d2, d3);
	nor (d7, d1);
	buf (d8, d2);
	or (d9, d2, d3);
	and (d10, d2, d4);
	xor (d11, d1, d4);
	not (d12, x1);
	and (d13, d1, d4);
	and (d14, d1);
	xor (d15, d1, d3);
	xor (d16, d4);
	or (d17, d2, d4);
	nand (d18, d2);
	and (d19, d1, d2);
	xnor (d20, d1, d4);
	and (d21, d4);
	xnor (d22, d1);
	buf (d23, d4);
	nand (d24, d4);
	nand (d25, d2, d3);
	and (d26, d3, d4);
	xor (d27, d1, d4);
	not (d28, d2);
	xnor (d29, d1, d3);
	xnor (d30, d1, d4);
	xor (d31, d2, d3);
	or (d32, d1, d3);
	xnor (d33, d2, d4);
	xor (d34, d1, d3);
	or (d35, d1, d2);
	xor (d36, d3, d4);
	nand (d37, d18, d31);
	buf (d38, d8);
	xor (d39, d28, d32);
	and (d40, d29, d33);
	nor (d41, d22, d28);
	not (d42, d32);
	nand (d43, d11, d30);
	nor (d44, d9, d33);
	buf (d45, d3);
	buf (d46, d25);
	and (d47, d8, d14);
	buf (d48, d35);
	or (d49, d11, d33);
	or (d50, d8, d33);
	xor (d51, d32, d36);
	nand (d52, d12, d32);
	nand (d53, d12, d16);
	and (d54, d28, d32);
	xor (d55, d13, d35);
	nor (d56, d9, d36);
	and (d57, d27, d31);
	or (d58, d10, d36);
	nor (d59, d12, d31);
	nand (d60, d38, d48);
	not (d61, d40);
	nand (d62, d45, d57);
	xor (d63, d42, d55);
	or (d64, d52, d57);
	nor (d65, d37, d50);
	buf (d66, d9);
	nor (d67, d47, d54);
	xor (d68, d39, d41);
	and (d69, d37, d48);
	xnor (d70, d43, d58);
	and (d71, d48, d58);
	not (d72, d3);
	buf (d73, d32);
	and (d74, d41, d43);
	not (d75, d17);
	nand (d76, d39, d44);
	or (d77, d59);
	xor (d78, d43, d55);
	not (d79, d35);
	or (d80, d46, d59);
	buf (d81, d47);
	not (d82, d39);
	xor (d83, d43, d49);
	buf (d84, d41);
	xnor (d85, d43, d55);
	and (d86, d40, d41);
	not (d87, d58);
	nor (d88, d37, d53);
	xnor (d89, d49, d56);
	xor (d90, d38, d46);
	or (d91, d41, d55);
	nor (d92, d49);
	not (d93, d49);
	or (d94, d38, d50);
	nor (d95, d48, d49);
	or (d96, d43, d56);
	xor (d97, d46, d48);
	nor (d98, d37, d55);
	and (d99, d39, d57);
	not (d100, d25);
	nand (d101, d42, d45);
	nand (d102, d54, d57);
	and (d103, d45, d48);
	and (d104, d37, d51);
	or (d105, d39, d55);
	or (d106, d39, d56);
	xnor (d107, d41, d53);
	not (d108, d4);
	xor (d109, d38, d54);
	or (d110, d41, d58);
	nor (d111, d43);
	xor (d112, d54, d55);
	nand (d113, d41, d57);
	xor (d114, d51, d59);
	not (d115, d18);
	or (d116, d47, d49);
	xor (d117, d38, d41);
	nand (d118, d39, d41);
	or (d119, d45, d47);
	buf (d120, d42);
	and (d121, d39, d58);
	or (d122, d52, d55);
	nand (d123, d47, d57);
	not (d124, d30);
	not (d125, d27);
	nand (d126, d45, d49);
	nor (d127, d57, d59);
	not (d128, d8);
	xor (d129, d47, d57);
	xor (d130, d50, d58);
	not (d131, d44);
	not (d132, d21);
	nand (d133, d50, d51);
	nand (d134, d45);
	nand (d135, d47, d59);
	nor (d136, d45, d52);
	nor (d137, d38, d58);
	nand (d138, d37, d49);
	nand (d139, d39, d50);
	xor (d140, d55, d59);
	nand (d141, d56, d59);
	xnor (d142, d46, d56);
	not (d143, d10);
	assign f1 = d60;
	assign f2 = d118;
	assign f3 = d80;
	assign f4 = d66;
	assign f5 = d81;
endmodule
