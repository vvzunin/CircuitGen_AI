module CCGRCG190( x0, x1, x2, x3, x4, x5, x6, f1, f2 );

	input x0, x1, x2, x3, x4, x5, x6;
	output f1, f2;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292;

	nand (d1, x1, x6);
	or (d2, x2, x5);
	xor (d3, x1, x4);
	xnor (d4, x2, x6);
	xnor (d5, x0, x6);
	and (d6, x3);
	and (d7, x2, x4);
	and (d8, x3, x6);
	nor (d9, x1, x6);
	nor (d10, x3, x4);
	xor (d11, x3, x6);
	buf (d12, x1);
	nand (d13, x4);
	nor (d14, x0, x1);
	buf (d15, x5);
	and (d16, x6);
	or (d17, x6);
	and (d18, x0);
	buf (d19, x6);
	nand (d20, x0, x3);
	not (d21, x2);
	xor (d22, x0, x6);
	nand (d23, x6);
	not (d24, x0);
	xnor (d25, x0, x5);
	xor (d26, x2, x5);
	not (d27, x1);
	nand (d28, x3, x5);
	xnor (d29, x2, x4);
	or (d30, x4, x5);
	buf (d31, x3);
	xor (d32, x4, x6);
	nand (d33, x0, x2);
	xor (d34, x0, x3);
	not (d35, x4);
	and (d36, x1, x3);
	nor (d37, x5, x6);
	buf (d38, x4);
	nor (d39, x4, x6);
	xnor (d40, x3, x4);
	nand (d41, x2, x5);
	or (d42, x1, x6);
	nor (d43, x1, x3);
	or (d44, x2, x5);
	and (d45, x2, x6);
	and (d46, x3, x4);
	xnor (d47, x0, x2);
	and (d48, x0, x2);
	nor (d49, x5, x6);
	nand (d50, x2, x5);
	and (d51, x5, x6);
	or (d52, x2, x3);
	xnor (d53, x1, x5);
	not (d54, x5);
	or (d55, x3, x5);
	xnor (d56, x0, x1);
	xnor (d57, x2, x3);
	xor (d58, x3);
	xor (d59, x5, x6);
	or (d60, x5);
	nand (d61, x5, x6);
	nand (d62, x2, x6);
	and (d63, x1, x5);
	nand (d64, x2, x4);
	or (d65, x3, x5);
	xor (d66, x3, x4);
	xor (d67, x2, x6);
	buf (d68, x2);
	xor (d69, x4, x6);
	xor (d70, x2, x4);
	not (d71, x3);
	xor (d72, x1, x2);
	or (d73, x4);
	xor (d74, x1);
	nor (d75, x3, x6);
	nor (d76, x1);
	nor (d77, x3, x4);
	and (d78, x1, x5);
	xor (d79, x2);
	buf (d80, d13);
	not (d81, d54);
	or (d82, d48, d55);
	and (d83, d69, d78);
	or (d84, d7, d77);
	or (d85, d10, d42);
	xnor (d86, d59, d67);
	nand (d87, d32, d78);
	nor (d88, d15, d49);
	and (d89, d58, d72);
	and (d90, d11, d63);
	and (d91, d2, d28);
	not (d92, d71);
	or (d93, d2, d58);
	xnor (d94, d13, d71);
	nor (d95, d55, d63);
	not (d96, d46);
	or (d97, d20, d55);
	buf (d98, d19);
	nor (d99, d31, d61);
	xor (d100, d24, d58);
	or (d101, d61, d64);
	nand (d102, d28, d76);
	xor (d103, d8, d40);
	and (d104, d60, d76);
	xnor (d105, d2, d14);
	or (d106, d39, d43);
	or (d107, d2, d31);
	xnor (d108, d45, d56);
	or (d109, d27, d35);
	nand (d110, d53, d60);
	nand (d111, d21, d57);
	not (d112, d4);
	buf (d113, d79);
	nor (d114, d6, d36);
	not (d115, d42);
	nand (d116, d2, d19);
	buf (d117, d63);
	nor (d118, d7, d69);
	buf (d119, d1);
	xnor (d120, d7, d62);
	not (d121, d19);
	xor (d122, d2, d3);
	not (d123, d57);
	xor (d124, d33, d71);
	or (d125, d27, d79);
	and (d126, d60, d63);
	and (d127, d12, d59);
	and (d128, d3, d69);
	buf (d129, d47);
	nand (d130, d50, d54);
	buf (d131, d4);
	xnor (d132, d10, d62);
	and (d133, d12, d25);
	xor (d134, d34, d62);
	or (d135, d7, d33);
	not (d136, d52);
	xnor (d137, d12, d24);
	nor (d138, d32, d77);
	nand (d139, d71, d72);
	and (d140, d15, d75);
	buf (d141, d32);
	nor (d142, d18, d64);
	buf (d143, d75);
	and (d144, d34, d36);
	nand (d145, d19, d41);
	buf (d146, d60);
	nor (d147, d47, d78);
	and (d148, d11, d49);
	and (d149, d108, d125);
	and (d150, d139, d148);
	nand (d151, d95, d142);
	nor (d152, d86, d87);
	buf (d153, d93);
	nor (d154, d124, d143);
	xnor (d155, d97, d122);
	and (d156, d103, d144);
	nor (d157, d105, d146);
	not (d158, d38);
	xnor (d159, d112, d142);
	xnor (d160, d91, d108);
	or (d161, d131, d146);
	xnor (d162, d142, d147);
	nand (d163, d92, d114);
	and (d164, d80, d117);
	nor (d165, d85, d101);
	xnor (d166, d82, d99);
	or (d167, d91, d128);
	xor (d168, d105, d139);
	not (d169, d56);
	not (d170, d60);
	nor (d171, d126, d146);
	or (d172, d115, d132);
	nor (d173, d97, d128);
	not (d174, d102);
	or (d175, d121, d135);
	buf (d176, d147);
	nand (d177, d82, d121);
	buf (d178, d27);
	xnor (d179, d119, d139);
	or (d180, d109);
	and (d181, d81, d101);
	nor (d182, d90, d96);
	or (d183, d122, d146);
	xnor (d184, d120, d131);
	xnor (d185, d90, d147);
	nand (d186, d86, d90);
	and (d187, d119, d148);
	buf (d188, d33);
	buf (d189, d121);
	xnor (d190, d84, d98);
	nor (d191, d83, d86);
	and (d192, d108, d141);
	buf (d193, d117);
	buf (d194, d21);
	nand (d195, d119, d147);
	or (d196, d120, d135);
	xnor (d197, d117, d131);
	nor (d198, d89, d147);
	xnor (d199, d89, d98);
	nor (d200, d86, d126);
	nor (d201, d87, d97);
	nand (d202, d93, d119);
	not (d203, d58);
	xnor (d204, d166, d185);
	xor (d205, d170, d197);
	xor (d206, d185, d195);
	not (d207, d132);
	buf (d208, d81);
	nand (d209, d191, d197);
	and (d210, d157, d161);
	or (d211, d154, d199);
	or (d212, d150, d171);
	not (d213, d175);
	not (d214, d167);
	nand (d215, d149, d190);
	xnor (d216, d161, d179);
	nor (d217, d162, d190);
	and (d218, d154, d182);
	buf (d219, d154);
	and (d220, d151, d174);
	nand (d221, d171, d194);
	and (d222, d160, d168);
	xnor (d223, d155, d200);
	nand (d224, d181, d187);
	not (d225, d25);
	nor (d226, d152, d161);
	nand (d227, d176, d198);
	nor (d228, d151, d179);
	not (d229, d186);
	xor (d230, d163, d187);
	nand (d231, d150, d183);
	or (d232, d151, d170);
	xor (d233, d174, d177);
	or (d234, d162, d200);
	nand (d235, d176, d183);
	buf (d236, d51);
	nor (d237, d184, d193);
	nand (d238, d156, d168);
	not (d239, d77);
	nor (d240, d151, d188);
	nor (d241, d162, d186);
	not (d242, d44);
	buf (d243, d44);
	nor (d244, d162, d198);
	or (d245, d156, d165);
	buf (d246, d144);
	not (d247, d63);
	xor (d248, d163, d164);
	buf (d249, d30);
	nand (d250, d155, d169);
	nor (d251, d170, d187);
	not (d252, d172);
	buf (d253, d17);
	xor (d254, d150, d197);
	buf (d255, d72);
	nand (d256, d154, d161);
	not (d257, d135);
	nand (d258, d181, d191);
	or (d259, d149, d162);
	not (d260, d104);
	nand (d261, d152, d195);
	and (d262, d190, d192);
	xnor (d263, d150, d159);
	buf (d264, d95);
	buf (d265, d114);
	nand (d266, d153, d180);
	nand (d267, d183, d199);
	and (d268, d186, d192);
	xor (d269, d168, d189);
	or (d270, d154, d195);
	nand (d271, d154, d158);
	xor (d272, d176, d191);
	buf (d273, d125);
	nor (d274, d175, d195);
	xnor (d275, d170, d173);
	buf (d276, d139);
	xnor (d277, d173, d193);
	xnor (d278, d159, d181);
	not (d279, d100);
	or (d280, d170, d183);
	not (d281, d68);
	nand (d282, d158, d190);
	buf (d283, d122);
	and (d284, d152, d187);
	nor (d285, d177, d182);
	buf (d286, d175);
	not (d287, d128);
	or (d288, d178, d189);
	buf (d289, d68);
	nand (d290, d161, d195);
	or (d291, d163, d177);
	xor (d292, d164, d188);
	assign f1 = d214;
	assign f2 = d288;
endmodule
