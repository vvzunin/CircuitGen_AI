module CCGRCG105( x0, x1, x2, x3, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16 );

	input x0, x1, x2, x3;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237;

	buf (d1, x1);
	nor (d2, x0, x3);
	or (d3, x0, x3);
	buf (d4, x0);
	nor (d5, x1);
	xor (d6, x2, x3);
	xnor (d7, x1, x2);
	and (d8, x1, x2);
	nor (d9, x1, x2);
	xor (d10, x2);
	xnor (d11, x2, x3);
	xnor (d12, x1, x3);
	and (d13, x0, x1);
	or (d14, x0, x1);
	and (d15, x0, x3);
	not (d16, x1);
	or (d17, x0, x1);
	and (d18, x2, x3);
	and (d19, x1, x3);
	xor (d20, x1, x3);
	not (d21, x0);
	and (d22, x1, x3);
	nand (d23, x0, x3);
	xnor (d24, x0, x1);
	buf (d25, x2);
	or (d26, d6, d12);
	and (d27, d4, d20);
	nor (d28, d26);
	not (d29, d16);
	buf (d30, d26);
	xnor (d31, d26, d27);
	buf (d32, x3);
	or (d33, d27);
	nand (d34, d29, d31);
	xor (d35, d29, d32);
	xor (d36, d29);
	buf (d37, d16);
	nor (d38, d28, d32);
	xnor (d39, d31, d33);
	nor (d40, d31, d32);
	or (d41, d30, d33);
	xnor (d42, d28, d32);
	xor (d43, d31, d33);
	or (d44, d29, d30);
	xnor (d45, d33);
	xnor (d46, d30, d32);
	nand (d47, d28, d30);
	or (d48, d31, d32);
	not (d49, d13);
	nand (d50, d29, d30);
	not (d51, d11);
	buf (d52, d5);
	xor (d53, d28, d31);
	not (d54, x3);
	xor (d55, d28);
	not (d56, d14);
	xnor (d57, d32);
	buf (d58, d12);
	and (d59, d32, d33);
	xnor (d60, d31);
	xnor (d61, d28, d33);
	nand (d62, d29, d32);
	nor (d63, d59, d61);
	or (d64, d36, d57);
	or (d65, d35, d61);
	xor (d66, d36, d52);
	and (d67, d47, d53);
	not (d68, d18);
	not (d69, d21);
	nor (d70, d34, d44);
	xnor (d71, d64, d66);
	not (d72, d68);
	buf (d73, d68);
	xnor (d74, d66, d67);
	xor (d75, d63, d64);
	not (d76, d23);
	buf (d77, d67);
	buf (d78, d7);
	and (d79, d63, d67);
	buf (d80, d66);
	and (d81, d75, d79);
	and (d82, d73, d78);
	nand (d83, d72, d77);
	xnor (d84, d76, d79);
	xnor (d85, d72, d78);
	or (d86, d73, d74);
	and (d87, d74, d78);
	or (d88, d72);
	nor (d89, d74, d76);
	xor (d90, d75, d80);
	not (d91, d44);
	or (d92, d73, d75);
	xnor (d93, d77, d80);
	nand (d94, d73, d74);
	and (d95, d71, d75);
	or (d96, d76, d79);
	xnor (d97, d76, d78);
	xnor (d98, d73, d75);
	nor (d99, d78, d80);
	and (d100, d72, d73);
	xnor (d101, d75, d80);
	nor (d102, d77, d80);
	xnor (d103, d75, d77);
	or (d104, d72, d78);
	nor (d105, d72, d75);
	not (d106, d66);
	or (d107, d73, d74);
	and (d108, d71, d73);
	xor (d109, d72, d77);
	xnor (d110, d96, d102);
	nand (d111, d88, d98);
	buf (d112, d46);
	and (d113, d85, d86);
	xnor (d114, d98, d104);
	nand (d115, d85, d106);
	not (d116, d54);
	xor (d117, d101, d107);
	nor (d118, d101, d104);
	nand (d119, d103, d107);
	not (d120, d77);
	not (d121, d71);
	xor (d122, d99, d107);
	nor (d123, d85, d104);
	xor (d124, d86, d104);
	nand (d125, d93, d107);
	xor (d126, d85, d106);
	nand (d127, d89, d105);
	xnor (d128, d94);
	xor (d129, d94, d109);
	or (d130, d88, d107);
	buf (d131, d94);
	not (d132, d52);
	nand (d133, d102, d106);
	buf (d134, d10);
	or (d135, d103, d104);
	nor (d136, d125, d126);
	or (d137, d113, d124);
	xor (d138, d119, d126);
	buf (d139, d77);
	buf (d140, d18);
	buf (d141, d75);
	and (d142, d117, d128);
	nand (d143, d125);
	and (d144, d121, d134);
	not (d145, d104);
	nor (d146, d114, d131);
	xor (d147, d131);
	xor (d148, d113, d125);
	buf (d149, d121);
	buf (d150, d6);
	nand (d151, d111, d123);
	nand (d152, d131);
	not (d153, d25);
	or (d154, d115, d134);
	buf (d155, d134);
	nand (d156, d122, d131);
	nor (d157, d116, d132);
	nand (d158, d124, d128);
	buf (d159, d127);
	nand (d160, d118, d129);
	or (d161, d114, d123);
	nand (d162, d115, d128);
	and (d163, d115, d131);
	xor (d164, d111, d115);
	nor (d165, d117, d118);
	or (d166, d127, d129);
	and (d167, d117, d118);
	and (d168, d121, d132);
	not (d169, d37);
	xor (d170, d126, d131);
	or (d171, d110, d127);
	xor (d172, d117, d120);
	not (d173, d118);
	nand (d174, d125, d132);
	nand (d175, d112, d124);
	xor (d176, d125, d133);
	or (d177, d110, d132);
	nand (d178, d119, d124);
	or (d179, d127, d129);
	xnor (d180, d118, d130);
	nand (d181, d110, d117);
	xnor (d182, d110, d133);
	or (d183, d124, d126);
	xnor (d184, d118, d119);
	buf (d185, d29);
	buf (d186, d24);
	nor (d187, d121, d132);
	buf (d188, d123);
	buf (d189, d39);
	or (d190, d115, d120);
	and (d191, d150, d157);
	xnor (d192, d163);
	nand (d193, d145, d169);
	or (d194, d141, d147);
	and (d195, d162, d186);
	not (d196, d32);
	xor (d197, d172, d187);
	not (d198, d139);
	nand (d199, d146, d149);
	or (d200, d179, d185);
	nor (d201, d161, d168);
	nand (d202, d154, d178);
	xnor (d203, d163, d168);
	and (d204, d152, d164);
	not (d205, d8);
	xor (d206, d144, d158);
	buf (d207, d30);
	xnor (d208, d159, d182);
	buf (d209, d95);
	nor (d210, d154, d166);
	nand (d211, d161, d185);
	xor (d212, d150, d161);
	nor (d213, d136, d184);
	xnor (d214, d159, d173);
	or (d215, d175, d177);
	not (d216, d67);
	nor (d217, d146, d174);
	xor (d218, d180, d186);
	or (d219, d154, d181);
	xnor (d220, d144, d175);
	xnor (d221, d150, d173);
	xor (d222, d172, d180);
	and (d223, d170, d181);
	xnor (d224, d152, d153);
	not (d225, d186);
	buf (d226, d130);
	buf (d227, d88);
	xor (d228, d167, d168);
	and (d229, d144, d162);
	and (d230, d164, d180);
	xnor (d231, d158, d168);
	xor (d232, d153, d176);
	xor (d233, d172, d183);
	or (d234, d141, d161);
	not (d235, d70);
	and (d236, d144, d155);
	xnor (d237, d163, d181);
	assign f1 = d211;
	assign f2 = d193;
	assign f3 = d225;
	assign f4 = d222;
	assign f5 = d208;
	assign f6 = d221;
	assign f7 = d225;
	assign f8 = d218;
	assign f9 = d194;
	assign f10 = d231;
	assign f11 = d198;
	assign f12 = d203;
	assign f13 = d234;
	assign f14 = d216;
	assign f15 = d192;
	assign f16 = d217;
endmodule
