module CCGRCG111( x0, x1, x2, x3, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17, f18, f19 );

	input x0, x1, x2, x3;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17, f18, f19;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58;

	xnor (d1, x0, x3);
	buf (d2, x1);
	nand (d3, x1, x3);
	xor (d4, x0, x3);
	not (d5, x3);
	nand (d6, x2, x3);
	nor (d7, x0, x3);
	nand (d8, x2, x3);
	xnor (d9, x0, x2);
	xor (d10, x1, x3);
	nand (d11, x1, x2);
	and (d12, x3);
	buf (d13, x0);
	or (d14, x0, x1);
	xnor (d15, x2, x3);
	and (d16, x1, x2);
	and (d17, x0, x2);
	xnor (d18, x1, x2);
	xor (d19, x2, x3);
	and (d20, x1, x3);
	and (d21, x1, x3);
	nand (d22, x0, x1);
	or (d23, x2);
	buf (d24, x3);
	and (d25, x0, x1);
	nor (d26, x1, x2);
	nor (d27, x0, x1);
	or (d28, x3);
	xnor (d29, x0, x3);
	or (d30, x0, x2);
	or (d31, x0, x3);
	and (d32, x0, x2);
	and (d33, x2);
	or (d34, x1, x2);
	xor (d35, x1);
	nand (d36, x1, x2);
	nor (d37, x0, x2);
	not (d38, x2);
	or (d39, x1, x3);
	not (d40, x0);
	nand (d41, x0, x1);
	and (d42, x0, x3);
	or (d43, x0, x3);
	not (d44, x1);
	and (d45, x0, x3);
	nor (d46, x2);
	nor (d47, x2, x3);
	nand (d48, x1, x3);
	and (d49, x0, x1);
	nor (d50, x0);
	xor (d51, x0, x2);
	xnor (d52, x1, x2);
	xnor (d53, x2);
	or (d54, x0, x1);
	xor (d55, x2);
	and (d56, x0);
	xnor (d57, x0, x2);
	nor (d58, x1);
	assign f1 = d17;
	assign f2 = d14;
	assign f3 = d51;
	assign f4 = d3;
	assign f5 = d53;
	assign f6 = d47;
	assign f7 = d7;
	assign f8 = d3;
	assign f9 = d13;
	assign f10 = d32;
	assign f11 = d10;
	assign f12 = d30;
	assign f13 = d1;
	assign f14 = d12;
	assign f15 = d14;
	assign f16 = d53;
	assign f17 = d48;
	assign f18 = d7;
	assign f19 = d16;
endmodule
