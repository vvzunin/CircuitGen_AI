module CCGRCG7( x0, x1, f1, f2, f3, f4, f5 );

	input x0, x1;
	output f1, f2, f3, f4, f5;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314, d315, d316, d317, d318, d319, d320, d321, d322, d323, d324, d325, d326, d327, d328, d329, d330, d331, d332, d333, d334, d335, d336, d337, d338, d339, d340, d341, d342, d343, d344, d345, d346, d347, d348, d349, d350, d351, d352, d353, d354, d355, d356, d357, d358, d359, d360, d361, d362, d363, d364, d365, d366, d367, d368, d369, d370;

	or (d1, x0, x1);
	buf (d2, x1);
	xor (d3, x0);
	nand (d4, x0, x1);
	xor (d5, x0, x1);
	not (d6, x0);
	xnor (d7, x1);
	nand (d8, x0, x1);
	nand (d9, x0);
	xor (d10, x1);
	or (d11, x0, x1);
	buf (d12, x0);
	and (d13, x0);
	nor (d14, x0);
	and (d15, x0, x1);
	and (d16, x0, x1);
	xnor (d17, x0, x1);
	xnor (d18, x0);
	not (d19, x1);
	or (d20, x1);
	xnor (d21, x0, x1);
	nand (d22, x1);
	or (d23, x0);
	xor (d24, x0, x1);
	nor (d25, x0, x1);
	xor (d26, d12, d25);
	nand (d27, d16, d22);
	or (d28, d5, d23);
	and (d29, d10, d16);
	nand (d30, d10, d22);
	nor (d31, d8, d15);
	nand (d32, d19, d22);
	xnor (d33, d6, d22);
	nor (d34, d16, d17);
	not (d35, d20);
	not (d36, d5);
	or (d37, d3, d13);
	nand (d38, d10, d11);
	or (d39, d21, d24);
	or (d40, d6, d8);
	buf (d41, d17);
	and (d42, d11, d20);
	or (d43, d4, d23);
	xnor (d44, d18, d24);
	nand (d45, d7, d19);
	buf (d46, d8);
	xnor (d47, d9, d21);
	or (d48, d1, d16);
	and (d49, d10, d21);
	nand (d50, d20, d22);
	and (d51, d1, d13);
	not (d52, d17);
	nand (d53, d9, d13);
	nor (d54, d2, d8);
	xor (d55, d25);
	xor (d56, d12, d13);
	or (d57, d3, d21);
	nand (d58, d14, d20);
	xnor (d59, d5, d8);
	xor (d60, d4, d20);
	buf (d61, d20);
	or (d62, d5, d21);
	xnor (d63, d11, d21);
	not (d64, d15);
	or (d65, d22, d25);
	nor (d66, d13, d15);
	nor (d67, d19, d25);
	buf (d68, d19);
	or (d69, d5, d8);
	nor (d70, d3, d6);
	xor (d71, d1, d21);
	xnor (d72, d24, d25);
	not (d73, d18);
	not (d74, d8);
	nor (d75, d2, d11);
	xor (d76, d30, d44);
	and (d77, d45, d75);
	nor (d78, d48, d51);
	xnor (d79, d54, d71);
	xnor (d80, d38, d69);
	nand (d81, d40, d72);
	and (d82, d29, d40);
	nor (d83, d38, d63);
	xnor (d84, d64, d67);
	and (d85, d62, d72);
	xnor (d86, d43, d61);
	not (d87, d41);
	and (d88, d45, d54);
	nand (d89, d29, d42);
	nor (d90, d31, d48);
	xor (d91, d54, d75);
	or (d92, d35, d71);
	xnor (d93, d36, d55);
	xnor (d94, d45, d65);
	buf (d95, d14);
	buf (d96, d24);
	buf (d97, d42);
	xnor (d98, d64, d65);
	or (d99, d28, d32);
	xor (d100, d40, d53);
	xor (d101, d28, d53);
	and (d102, d36, d74);
	or (d103, d54, d60);
	nand (d104, d47, d66);
	not (d105, d14);
	nand (d106, d38, d73);
	nor (d107, d32, d51);
	and (d108, d28, d44);
	buf (d109, d32);
	and (d110, d27, d67);
	nor (d111, d27, d41);
	xnor (d112, d35, d38);
	or (d113, d37, d64);
	and (d114, d49);
	nor (d115, d34, d59);
	xor (d116, d36, d47);
	not (d117, d63);
	not (d118, d54);
	nand (d119, d55, d64);
	or (d120, d35, d63);
	or (d121, d35, d52);
	nor (d122, d28, d58);
	xnor (d123, d53, d57);
	and (d124, d33, d50);
	not (d125, d68);
	and (d126, d47, d54);
	nand (d127, d26, d48);
	nor (d128, d38, d48);
	not (d129, d57);
	nand (d130, d59, d66);
	nand (d131, d29, d70);
	not (d132, d47);
	buf (d133, d56);
	nor (d134, d55, d71);
	buf (d135, d69);
	nor (d136, d41, d75);
	nor (d137, d32, d33);
	xnor (d138, d67, d69);
	not (d139, d35);
	buf (d140, d49);
	not (d141, d26);
	xnor (d142, d32, d53);
	or (d143, d45, d48);
	xnor (d144, d36, d39);
	nand (d145, d29, d37);
	not (d146, d28);
	not (d147, d25);
	nand (d148, d112, d113);
	nand (d149, d84, d89);
	nand (d150, d124, d141);
	nand (d151, d111, d144);
	buf (d152, d77);
	or (d153, d137);
	xnor (d154, d102, d126);
	or (d155, d97, d126);
	xor (d156, d85, d140);
	nand (d157, d76, d136);
	and (d158, d134, d137);
	xnor (d159, d89, d117);
	and (d160, d83, d98);
	and (d161, d100, d122);
	xnor (d162, d94, d119);
	or (d163, d81, d135);
	nor (d164, d82, d131);
	buf (d165, d75);
	buf (d166, d143);
	buf (d167, d47);
	not (d168, d128);
	xnor (d169, d85, d90);
	nand (d170, d113, d130);
	xnor (d171, d132, d144);
	xor (d172, d113, d126);
	xnor (d173, d109, d114);
	buf (d174, d10);
	xor (d175, d80, d96);
	xnor (d176, d111, d116);
	not (d177, d1);
	xor (d178, d81, d85);
	and (d179, d102, d120);
	nor (d180, d82, d114);
	xnor (d181, d80, d128);
	not (d182, d121);
	xor (d183, d88, d145);
	buf (d184, d117);
	nand (d185, d77, d107);
	xor (d186, d130, d137);
	nand (d187, d88, d127);
	xor (d188, d129, d147);
	nor (d189, d87, d113);
	nor (d190, d82, d92);
	buf (d191, d44);
	buf (d192, d126);
	not (d193, d102);
	xnor (d194, d112, d137);
	xnor (d195, d108, d133);
	or (d196, d136, d138);
	and (d197, d79, d81);
	buf (d198, d142);
	xor (d199, d108, d127);
	nor (d200, d130);
	or (d201, d77, d96);
	xor (d202, d105, d132);
	xnor (d203, d128, d140);
	xor (d204, d79, d122);
	and (d205, d111, d118);
	nand (d206, d79, d119);
	buf (d207, d130);
	or (d208, d86, d98);
	buf (d209, d71);
	not (d210, d119);
	xor (d211, d77, d95);
	and (d212, d79, d138);
	not (d213, d13);
	not (d214, d78);
	nand (d215, d95, d142);
	or (d216, d88, d106);
	buf (d217, d96);
	xnor (d218, d114, d132);
	nand (d219, d93, d111);
	not (d220, d97);
	xnor (d221, d83, d115);
	xor (d222, d85, d128);
	xnor (d223, d89, d107);
	nand (d224, d108, d115);
	not (d225, d67);
	xor (d226, d114, d128);
	nand (d227, d94, d95);
	nor (d228, d88, d134);
	nand (d229, d91, d97);
	buf (d230, d114);
	buf (d231, d27);
	nor (d232, d119, d145);
	xor (d233, d95, d128);
	buf (d234, d128);
	buf (d235, d41);
	xor (d236, d95, d113);
	buf (d237, d36);
	nand (d238, d78, d92);
	xnor (d239, d114, d140);
	nor (d240, d118, d129);
	xnor (d241, d95, d147);
	buf (d242, d106);
	and (d243, d153, d219);
	and (d244, d177, d219);
	and (d245, d177, d217);
	nor (d246, d162, d165);
	and (d247, d206, d225);
	xor (d248, d204, d223);
	or (d249, d149, d156);
	buf (d250, d99);
	xnor (d251, d170, d176);
	or (d252, d149, d167);
	nand (d253, d151, d181);
	nor (d254, d150, d206);
	or (d255, d202, d210);
	nand (d256, d196, d199);
	nand (d257, d197, d241);
	or (d258, d188, d213);
	nor (d259, d209, d225);
	not (d260, d61);
	xnor (d261, d197, d204);
	nand (d262, d215, d234);
	nand (d263, d181, d215);
	or (d264, d195, d214);
	xnor (d265, d179, d229);
	nand (d266, d166, d181);
	buf (d267, d116);
	and (d268, d192, d204);
	xnor (d269, d217, d233);
	buf (d270, d132);
	xor (d271, d179, d228);
	and (d272, d150, d236);
	and (d273, d205, d234);
	xor (d274, d152, d193);
	xnor (d275, d154, d210);
	xor (d276, d214, d241);
	or (d277, d162, d168);
	xnor (d278, d171, d236);
	nor (d279, d195, d227);
	not (d280, d87);
	xor (d281, d268, d269);
	nand (d282, d254, d270);
	nor (d283, d265, d270);
	not (d284, d160);
	or (d285, d274, d278);
	or (d286, d242, d248);
	nor (d287, d250, d255);
	or (d288, d276, d279);
	nand (d289, d243, d277);
	or (d290, d270, d274);
	xnor (d291, d279);
	nand (d292, d242, d279);
	and (d293, d245, d266);
	and (d294, d258, d263);
	xnor (d295, d246, d249);
	nand (d296, d243, d262);
	nor (d297, d256, d261);
	or (d298, d251, d256);
	buf (d299, d3);
	or (d300, d267, d274);
	not (d301, d256);
	and (d302, d242, d247);
	xor (d303, d248, d262);
	nor (d304, d254, d259);
	xor (d305, d254, d265);
	and (d306, d245, d275);
	or (d307, d242, d277);
	xnor (d308, d270, d276);
	buf (d309, d273);
	and (d310, d243, d263);
	nand (d311, d260, d264);
	xnor (d312, d263, d264);
	xnor (d313, d270, d279);
	xor (d314, d243, d267);
	or (d315, d250, d259);
	or (d316, d247);
	xnor (d317, d272, d276);
	not (d318, d44);
	xor (d319, d263, d269);
	nand (d320, d249, d254);
	and (d321, d266);
	nor (d322, d265, d266);
	not (d323, d16);
	or (d324, d245, d268);
	xor (d325, d249, d251);
	nand (d326, d270, d272);
	xnor (d327, d245, d258);
	buf (d328, d84);
	nand (d329, d244, d246);
	not (d330, d221);
	xor (d331, d245, d259);
	and (d332, d275, d279);
	xnor (d333, d253, d268);
	xor (d334, d257, d265);
	nand (d335, d245, d262);
	nor (d336, d253, d272);
	xor (d337, d244, d272);
	nand (d338, d262, d275);
	xnor (d339, d261, d270);
	nand (d340, d249, d264);
	nand (d341, d244, d249);
	buf (d342, d129);
	xnor (d343, d248, d279);
	buf (d344, d67);
	xnor (d345, d266, d271);
	xor (d346, d247, d267);
	and (d347, d243, d257);
	nor (d348, d254, d270);
	nand (d349, d259, d270);
	xor (d350, d254, d267);
	not (d351, d9);
	xor (d352, d264, d278);
	nor (d353, d249, d278);
	nor (d354, d244, d262);
	nor (d355, d247, d262);
	buf (d356, d242);
	and (d357, d242, d273);
	and (d358, d258, d273);
	and (d359, d252, d263);
	nor (d360, d254, d277);
	buf (d361, d46);
	xnor (d362, d256, d265);
	or (d363, d249, d260);
	buf (d364, d185);
	and (d365, d264, d274);
	xor (d366, d244, d263);
	nand (d367, d270, d276);
	nor (d368, d256, d275);
	xor (d369, d261, d269);
	nor (d370, d242, d250);
	assign f1 = d307;
	assign f2 = d345;
	assign f3 = d338;
	assign f4 = d302;
	assign f5 = d336;
endmodule
