module CCGRCG89( x0, x1, x2, x3, f1, f2, f3, f4, f5, f6, f7, f8 );

	input x0, x1, x2, x3;
	output f1, f2, f3, f4, f5, f6, f7, f8;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314, d315, d316, d317, d318, d319, d320, d321, d322, d323, d324, d325, d326, d327, d328, d329, d330, d331, d332, d333, d334, d335, d336, d337, d338, d339, d340, d341, d342, d343, d344, d345, d346, d347, d348, d349, d350, d351, d352, d353, d354, d355, d356, d357, d358, d359, d360, d361, d362, d363, d364, d365, d366, d367, d368, d369, d370, d371, d372, d373, d374, d375, d376, d377, d378, d379, d380, d381, d382, d383, d384, d385, d386, d387, d388, d389, d390, d391, d392, d393, d394, d395, d396, d397, d398, d399, d400, d401, d402, d403, d404, d405, d406, d407, d408, d409, d410, d411, d412, d413, d414, d415, d416, d417, d418, d419, d420, d421, d422, d423, d424, d425, d426, d427, d428, d429, d430, d431, d432, d433, d434, d435, d436, d437, d438, d439, d440, d441, d442, d443, d444, d445, d446, d447, d448, d449, d450, d451, d452, d453, d454, d455, d456, d457, d458, d459, d460, d461, d462, d463, d464;

	nand (d1, x1, x3);
	buf (d2, x1);
	not (d3, x1);
	nand (d4, x0);
	nor (d5, x3);
	nand (d6, x0, x2);
	nor (d7, x0);
	xor (d8, x1, x2);
	xor (d9, x3);
	nor (d10, x2);
	xnor (d11, x1, x3);
	nor (d12, d1, d7);
	nor (d13, d3, d9);
	buf (d14, d10);
	xor (d15, d3, d11);
	xnor (d16, d2, d10);
	nor (d17, d1, d5);
	and (d18, d7, d10);
	or (d19, d1, d8);
	xor (d20, d10);
	nor (d21, d6);
	nor (d22, d7, d8);
	xnor (d23, d7, d8);
	nor (d24, d8, d10);
	nand (d25, d7, d9);
	buf (d26, d4);
	xor (d27, d3, d9);
	not (d28, d4);
	xnor (d29, d9, d11);
	nand (d30, d6, d7);
	and (d31, d3, d4);
	nor (d32, d5);
	xor (d33, d6, d10);
	xnor (d34, d8, d10);
	buf (d35, x2);
	buf (d36, d1);
	xor (d37, d10, d11);
	and (d38, d7, d9);
	and (d39, d4, d9);
	xnor (d40, d1, d5);
	not (d41, x2);
	nand (d42, d6, d8);
	not (d43, d2);
	not (d44, d11);
	or (d45, d2, d8);
	or (d46, d3, d8);
	or (d47, d1, d2);
	xnor (d48, d3, d4);
	nor (d49, d1, d7);
	nand (d50, d2, d6);
	xor (d51, d9, d11);
	buf (d52, d11);
	and (d53, d2);
	xor (d54, d5, d8);
	or (d55, d10, d11);
	xor (d56, d2, d10);
	or (d57, d3, d10);
	not (d58, x0);
	buf (d59, d8);
	or (d60, d2, d5);
	nor (d61, d4, d6);
	buf (d62, d3);
	xor (d63, d6, d7);
	nor (d64, d5, d8);
	nand (d65, d7);
	not (d66, d10);
	xnor (d67, d3, d6);
	xor (d68, d2, d10);
	xnor (d69, d6, d7);
	and (d70, d4, d6);
	xor (d71, d2, d5);
	nor (d72, d1, d6);
	xor (d73, d3, d7);
	xor (d74, d7, d9);
	xor (d75, d6, d9);
	xnor (d76, d9, d11);
	or (d77, d2);
	xnor (d78, d3, d7);
	not (d79, d8);
	nand (d80, d3, d9);
	buf (d81, d7);
	nor (d82, d4, d7);
	xnor (d83, d5, d10);
	or (d84, d6, d9);
	nand (d85, d31, d79);
	xor (d86, d18);
	and (d87, d22, d69);
	nand (d88, d16, d39);
	buf (d89, d29);
	xnor (d90, d56, d79);
	xnor (d91, d47, d54);
	xnor (d92, d35, d74);
	or (d93, d39, d40);
	nor (d94, d14, d81);
	nand (d95, d12, d83);
	or (d96, d33, d63);
	nand (d97, d50, d62);
	buf (d98, d83);
	xnor (d99, d51, d81);
	or (d100, d33, d78);
	and (d101, d91, d95);
	nor (d102, d93, d98);
	nand (d103, d86, d97);
	or (d104, d89, d95);
	nor (d105, d87, d97);
	nor (d106, d85, d98);
	nand (d107, d87, d100);
	xnor (d108, d89, d92);
	buf (d109, d33);
	and (d110, d99, d100);
	xor (d111, d87, d88);
	buf (d112, d42);
	buf (d113, d48);
	and (d114, d91, d93);
	nor (d115, d88, d99);
	xnor (d116, d86, d93);
	and (d117, d86, d93);
	xnor (d118, d85, d88);
	or (d119, d94, d100);
	xor (d120, d92, d93);
	nand (d121, d95, d96);
	nor (d122, d86, d87);
	xnor (d123, d85, d100);
	and (d124, d90, d95);
	or (d125, d85, d92);
	xnor (d126, d100);
	xnor (d127, d86, d87);
	not (d128, d99);
	nand (d129, d86, d99);
	and (d130, d91, d98);
	not (d131, d29);
	or (d132, d90, d100);
	and (d133, d88, d93);
	xor (d134, d90, d91);
	and (d135, d92, d99);
	buf (d136, d76);
	nor (d137, d93, d94);
	buf (d138, d91);
	xor (d139, d86, d95);
	and (d140, d92, d95);
	xor (d141, d86, d97);
	and (d142, d91, d94);
	xor (d143, d86, d100);
	nor (d144, d86, d92);
	xnor (d145, d96, d100);
	nand (d146, d96, d99);
	or (d147, d98, d100);
	not (d148, d42);
	not (d149, d36);
	or (d150, d85, d97);
	buf (d151, d84);
	xnor (d152, d92, d94);
	or (d153, d88, d97);
	xor (d154, d97, d100);
	xor (d155, d85, d100);
	xor (d156, d118, d126);
	xor (d157, d116, d123);
	xnor (d158, d133, d144);
	xor (d159, d112, d140);
	xnor (d160, d122, d129);
	and (d161, d108, d119);
	or (d162, d110, d128);
	nor (d163, d102, d117);
	nor (d164, d108, d110);
	nor (d165, d128, d155);
	not (d166, d101);
	xor (d167, d141, d152);
	or (d168, d128, d155);
	or (d169, d112, d117);
	or (d170, d108, d130);
	nor (d171, d122, d126);
	xnor (d172, d144, d148);
	and (d173, d139);
	not (d174, d78);
	not (d175, d135);
	and (d176, d114, d142);
	buf (d177, d5);
	or (d178, d110, d152);
	xor (d179, d113, d127);
	not (d180, d57);
	and (d181, d109, d143);
	not (d182, d65);
	not (d183, d71);
	or (d184, d121, d139);
	buf (d185, d147);
	nand (d186, d110, d111);
	buf (d187, d107);
	and (d188, d118, d130);
	not (d189, d147);
	nand (d190, d129, d136);
	xor (d191, d125, d149);
	and (d192, d129, d153);
	xnor (d193, d102, d137);
	not (d194, d70);
	xnor (d195, d110, d122);
	not (d196, d32);
	buf (d197, d80);
	nand (d198, d133, d136);
	xor (d199, d115, d148);
	or (d200, d116, d127);
	nand (d201, d125, d141);
	not (d202, d51);
	xnor (d203, d111, d152);
	nor (d204, d138, d152);
	nand (d205, d125, d134);
	xnor (d206, d101, d125);
	or (d207, d101, d154);
	or (d208, d130, d147);
	nor (d209, d115, d119);
	not (d210, d26);
	nor (d211, d135, d140);
	nor (d212, d109, d134);
	xnor (d213, d125, d152);
	or (d214, d105, d142);
	and (d215, d110, d147);
	and (d216, d104, d126);
	and (d217, d136, d152);
	xnor (d218, d105, d128);
	and (d219, d146, d152);
	nand (d220, d129, d150);
	xnor (d221, d102, d114);
	xnor (d222, d122, d127);
	xor (d223, d107, d147);
	xor (d224, d126, d147);
	and (d225, d103, d114);
	xnor (d226, d116, d155);
	nand (d227, d130, d144);
	xor (d228, d103, d150);
	not (d229, d48);
	nor (d230, d125, d141);
	xor (d231, d115, d125);
	and (d232, d115, d126);
	xnor (d233, d101, d146);
	xnor (d234, d101, d104);
	buf (d235, d68);
	xor (d236, d153, d154);
	or (d237, d104, d131);
	xnor (d238, d140, d144);
	or (d239, d119, d147);
	and (d240, d104, d152);
	buf (d241, d14);
	buf (d242, d122);
	xor (d243, d119, d130);
	buf (d244, d62);
	xnor (d245, d115, d144);
	nor (d246, d112, d117);
	nor (d247, d136, d155);
	not (d248, d130);
	or (d249, d106, d110);
	not (d250, d118);
	not (d251, d156);
	and (d252, d216, d238);
	nand (d253, d222, d248);
	not (d254, d201);
	nand (d255, d184, d214);
	buf (d256, d175);
	xor (d257, d171, d237);
	and (d258, d207, d241);
	and (d259, d156, d196);
	not (d260, d12);
	and (d261, d245, d249);
	xnor (d262, d167, d249);
	xnor (d263, d225, d231);
	and (d264, d177, d230);
	or (d265, d157, d203);
	or (d266, d170, d209);
	xor (d267, d181, d239);
	nand (d268, d198, d232);
	buf (d269, d235);
	and (d270, d209, d220);
	xnor (d271, d165, d230);
	and (d272, d174, d217);
	xnor (d273, d162, d208);
	nand (d274, d202, d242);
	nor (d275, d156, d206);
	or (d276, d200, d248);
	xor (d277, d163, d164);
	nand (d278, d201, d212);
	or (d279, d216, d227);
	xor (d280, d220, d230);
	xnor (d281, d205, d231);
	xnor (d282, d159, d242);
	xor (d283, d172, d183);
	or (d284, d196, d217);
	not (d285, d114);
	not (d286, d53);
	buf (d287, d150);
	buf (d288, d2);
	not (d289, d56);
	xor (d290, d166, d180);
	not (d291, x3);
	not (d292, d159);
	and (d293, d172, d246);
	buf (d294, d206);
	and (d295, d159, d210);
	or (d296, d175, d196);
	nand (d297, d227, d250);
	or (d298, d226, d228);
	and (d299, d159, d183);
	buf (d300, d226);
	xnor (d301, d225, d243);
	and (d302, d199, d222);
	or (d303, d165, d184);
	nor (d304, d173, d176);
	xnor (d305, d185, d222);
	xnor (d306, d172, d218);
	not (d307, d150);
	nand (d308, d167, d178);
	or (d309, d185, d201);
	xnor (d310, d223, d240);
	nand (d311, d189, d228);
	and (d312, d189, d243);
	xor (d313, d208, d225);
	xor (d314, d161, d245);
	xnor (d315, d181, d240);
	nor (d316, d183, d188);
	xnor (d317, d172, d191);
	xnor (d318, d173, d229);
	or (d319, d171, d238);
	xor (d320, d178, d220);
	xnor (d321, d174, d203);
	xnor (d322, d272, d321);
	and (d323, d286, d317);
	xor (d324, d256, d266);
	not (d325, d175);
	not (d326, d74);
	xnor (d327, d260, d310);
	nand (d328, d274, d277);
	buf (d329, d309);
	xnor (d330, d298, d305);
	not (d331, d191);
	and (d332, d269, d279);
	xnor (d333, d277, d302);
	nand (d334, d297, d319);
	buf (d335, d284);
	xnor (d336, d270, d296);
	nand (d337, d253, d320);
	xor (d338, d291, d301);
	nand (d339, d285, d310);
	xor (d340, d281, d317);
	nand (d341, d280, d314);
	nor (d342, d251, d259);
	xor (d343, d262, d276);
	nor (d344, d256, d260);
	and (d345, d262, d304);
	xor (d346, d266, d281);
	nand (d347, d268, d306);
	nor (d348, d291, d320);
	nand (d349, d265, d273);
	nand (d350, d269, d273);
	nor (d351, d273, d293);
	nand (d352, d295, d314);
	xnor (d353, d273, d294);
	nor (d354, d267, d279);
	and (d355, d282, d319);
	xor (d356, d272, d313);
	nor (d357, d251, d271);
	xnor (d358, d284, d296);
	and (d359, d281, d309);
	xor (d360, d272, d302);
	xnor (d361, d317, d319);
	buf (d362, d130);
	nand (d363, d263, d264);
	xnor (d364, d278, d321);
	xnor (d365, d290, d313);
	and (d366, d254, d272);
	xnor (d367, d270, d309);
	buf (d368, d124);
	nor (d369, d289, d296);
	xnor (d370, d268, d290);
	and (d371, d289, d300);
	or (d372, d252, d304);
	xor (d373, d276, d294);
	nand (d374, d299, d302);
	nand (d375, d263, d282);
	xor (d376, d253, d308);
	and (d377, d284, d312);
	not (d378, d186);
	and (d379, d313, d319);
	xnor (d380, d284, d321);
	nand (d381, d265, d307);
	and (d382, d270, d282);
	and (d383, d301, d305);
	not (d384, d161);
	nor (d385, d261, d287);
	buf (d386, d305);
	buf (d387, d69);
	or (d388, d288, d304);
	or (d389, d261, d266);
	not (d390, d47);
	not (d391, d293);
	not (d392, d239);
	buf (d393, d18);
	xnor (d394, d276, d292);
	and (d395, d298, d319);
	buf (d396, d58);
	nand (d397, d303, d310);
	nor (d398, d255, d295);
	buf (d399, d9);
	nand (d400, d283, d300);
	xor (d401, d296, d316);
	nor (d402, d257, d314);
	or (d403, d267, d291);
	not (d404, d52);
	and (d405, d285, d297);
	xor (d406, d322, d339);
	or (d407, d332, d338);
	xor (d408, d365, d396);
	not (d409, d391);
	nor (d410, d326, d341);
	buf (d411, d39);
	not (d412, d151);
	nor (d413, d388, d392);
	nand (d414, d335, d345);
	nor (d415, d348, d377);
	buf (d416, d44);
	buf (d417, d135);
	or (d418, d327, d359);
	nor (d419, d323, d336);
	xnor (d420, d362, d371);
	buf (d421, d263);
	nand (d422, d330, d398);
	xor (d423, d333, d399);
	not (d424, d103);
	xor (d425, d348, d398);
	xor (d426, d331, d332);
	nor (d427, d328, d383);
	or (d428, d395, d405);
	or (d429, d324, d349);
	xnor (d430, d379, d389);
	nor (d431, d361, d372);
	not (d432, d277);
	not (d433, d133);
	not (d434, d188);
	xor (d435, d369, d399);
	or (d436, d324, d365);
	xor (d437, d331, d396);
	or (d438, d338, d362);
	xor (d439, d350, d402);
	xnor (d440, d341, d376);
	nand (d441, d339, d388);
	nand (d442, d377, d384);
	buf (d443, d401);
	nand (d444, d387, d405);
	buf (d445, d174);
	xor (d446, d368, d383);
	or (d447, d330, d350);
	xnor (d448, d355, d377);
	or (d449, d369, d373);
	or (d450, d337, d354);
	not (d451, d30);
	xnor (d452, d359, d366);
	nor (d453, d335, d372);
	or (d454, d347, d401);
	nand (d455, d347, d385);
	or (d456, d323, d383);
	xor (d457, d324, d367);
	xnor (d458, d375, d398);
	xnor (d459, d355, d366);
	and (d460, d350, d381);
	buf (d461, d364);
	or (d462, d342, d385);
	buf (d463, d27);
	xnor (d464, d339, d360);
	assign f1 = d457;
	assign f2 = d432;
	assign f3 = d437;
	assign f4 = d462;
	assign f5 = d433;
	assign f6 = d437;
	assign f7 = d455;
	assign f8 = d437;
endmodule
