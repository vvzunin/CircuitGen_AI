module CCGRCG26( x0, x1, x2, f1, f2, f3, f4 );

	input x0, x1, x2;
	output f1, f2, f3, f4;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284;

	not (d1, x1);
	not (d2, x2);
	buf (d3, x1);
	buf (d4, x2);
	xnor (d5, x1);
	buf (d6, x0);
	xor (d7, x1, x2);
	nor (d8, x2);
	xor (d9, x2);
	not (d10, x0);
	and (d11, x0, x1);
	and (d12, x1);
	nand (d13, x0);
	xnor (d14, x0, x2);
	and (d15, x2);
	nand (d16, x1);
	or (d17, d6, d10);
	buf (d18, d7);
	xnor (d19, d4, d8);
	not (d20, d12);
	nand (d21, d13, d15);
	and (d22, d1, d3);
	nand (d23, d1, d11);
	nor (d24, d1, d11);
	xnor (d25, d5, d7);
	nor (d26, d8, d10);
	nor (d27, d21, d23);
	not (d28, d16);
	not (d29, d19);
	or (d30, d23, d26);
	nor (d31, d21, d26);
	nand (d32, d17, d24);
	xnor (d33, d21, d25);
	buf (d34, d12);
	not (d35, d18);
	not (d36, d4);
	and (d37, d24, d26);
	xor (d38, d19, d25);
	xor (d39, d20, d23);
	not (d40, d9);
	or (d41, d19, d24);
	nand (d42, d20, d24);
	buf (d43, d13);
	not (d44, d1);
	buf (d45, d22);
	xnor (d46, d30, d44);
	nand (d47, d41, d43);
	not (d48, d44);
	nor (d49, d36, d39);
	and (d50, d27, d33);
	nand (d51, d28, d37);
	xor (d52, d32, d40);
	nand (d53, d28, d34);
	or (d54, d42, d45);
	or (d55, d34, d36);
	xor (d56, d35, d37);
	not (d57, d35);
	and (d58, d38, d39);
	not (d59, d24);
	nor (d60, d28, d36);
	xor (d61, d29, d40);
	not (d62, d26);
	xnor (d63, d32, d35);
	nand (d64, d29, d32);
	or (d65, d36, d44);
	buf (d66, d38);
	not (d67, d13);
	xor (d68, d31, d36);
	not (d69, d34);
	and (d70, d31, d32);
	xnor (d71, d34, d45);
	xor (d72, d33, d37);
	or (d73, d33, d44);
	xnor (d74, d27, d35);
	nand (d75, d29, d36);
	xor (d76, d40, d45);
	and (d77, d29, d42);
	not (d78, d39);
	xnor (d79, d32, d38);
	or (d80, d29, d32);
	buf (d81, d1);
	not (d82, d15);
	or (d83, d27, d42);
	xor (d84, d38, d41);
	nor (d85, d31, d37);
	nand (d86, d27, d36);
	buf (d87, d41);
	or (d88, d41, d45);
	and (d89, d32, d45);
	buf (d90, d18);
	and (d91, d27, d33);
	nor (d92, d27, d33);
	nor (d93, d33, d38);
	xor (d94, d36, d44);
	nand (d95, d38, d45);
	nor (d96, d40, d43);
	nor (d97, d30, d44);
	and (d98, d29, d31);
	buf (d99, d40);
	or (d100, d33, d39);
	and (d101, d29, d37);
	buf (d102, d17);
	not (d103, d2);
	buf (d104, d26);
	nor (d105, d28, d45);
	xnor (d106, d43, d45);
	xor (d107, d31, d41);
	nor (d108, d28, d39);
	xnor (d109, d31, d33);
	xnor (d110, d31, d40);
	and (d111, d28, d32);
	nand (d112, d37, d45);
	or (d113, d33, d44);
	nor (d114, d36);
	and (d115, d30, d40);
	nor (d116, d39, d41);
	not (d117, d22);
	buf (d118, d39);
	nand (d119, d70, d84);
	nand (d120, d65, d66);
	or (d121, d102, d104);
	nand (d122, d61, d75);
	or (d123, d62, d83);
	xnor (d124, d93, d109);
	xnor (d125, d51, d56);
	xnor (d126, d85, d93);
	and (d127, d61, d106);
	nand (d128, d64, d95);
	and (d129, d57, d108);
	xnor (d130, d85, d97);
	nor (d131, d55, d72);
	buf (d132, d55);
	or (d133, d93, d116);
	not (d134, d114);
	and (d135, d76, d115);
	nor (d136, d101, d110);
	not (d137, d82);
	xnor (d138, d98, d107);
	and (d139, d50, d92);
	and (d140, d46, d55);
	or (d141, d69, d103);
	nor (d142, d74, d87);
	nor (d143, d57, d84);
	nand (d144, d62, d115);
	and (d145, d59, d90);
	or (d146, d91, d94);
	buf (d147, d10);
	or (d148, d119, d134);
	not (d149, d7);
	nand (d150, d126, d129);
	xnor (d151, d118, d137);
	not (d152, d41);
	and (d153, d139, d142);
	nor (d154, d128, d130);
	not (d155, d49);
	and (d156, d134, d140);
	xnor (d157, d124, d126);
	xor (d158, d136, d142);
	xnor (d159, d128, d131);
	nor (d160, d137, d146);
	xor (d161, d125, d138);
	nand (d162, d129, d141);
	buf (d163, d123);
	nand (d164, d118, d136);
	and (d165, d119, d142);
	nor (d166, d131, d136);
	or (d167, d128, d140);
	xnor (d168, d128, d135);
	xor (d169, d121, d141);
	buf (d170, d138);
	and (d171, d119, d125);
	nor (d172, d137, d144);
	xor (d173, d131, d143);
	nor (d174, d133, d140);
	xnor (d175, d138, d139);
	nor (d176, d123, d130);
	buf (d177, d101);
	or (d178, d128, d134);
	xor (d179, d138, d143);
	not (d180, d111);
	not (d181, d63);
	or (d182, d123, d132);
	nand (d183, d126, d130);
	or (d184, d129, d132);
	nor (d185, d129, d145);
	not (d186, d67);
	nor (d187, d126, d128);
	xor (d188, d123, d138);
	xor (d189, d125, d140);
	not (d190, d66);
	xnor (d191, d139, d142);
	and (d192, d121, d140);
	and (d193, d117, d140);
	and (d194, d130, d144);
	nor (d195, d119);
	not (d196, d77);
	not (d197, d102);
	xnor (d198, d129, d133);
	xnor (d199, d120, d146);
	xnor (d200, d119, d128);
	xnor (d201, d129);
	or (d202, d124, d125);
	or (d203, d120, d133);
	xor (d204, d143, d146);
	xor (d205, d142, d144);
	xor (d206, d132, d146);
	xnor (d207, d122, d141);
	buf (d208, d197);
	not (d209, d156);
	nand (d210, d158, d171);
	nand (d211, d168, d176);
	buf (d212, d92);
	and (d213, d150, d166);
	and (d214, d158, d175);
	xor (d215, d188, d199);
	and (d216, d152, d165);
	nand (d217, d162, d188);
	xnor (d218, d176, d182);
	buf (d219, d19);
	nor (d220, d184, d202);
	nor (d221, d182, d188);
	nor (d222, d190, d201);
	and (d223, d174, d197);
	nor (d224, d158, d195);
	nand (d225, d151, d180);
	or (d226, d162, d166);
	xor (d227, d181, d187);
	not (d228, d145);
	not (d229, d151);
	xor (d230, d186, d202);
	xnor (d231, d163, d205);
	and (d232, d152, d199);
	buf (d233, d180);
	and (d234, d151, d206);
	xnor (d235, d184, d200);
	nor (d236, d184, d186);
	nand (d237, d193, d206);
	buf (d238, d189);
	and (d239, d168, d203);
	and (d240, d194, d207);
	or (d241, d165, d189);
	xor (d242, d161, d167);
	xor (d243, d155, d191);
	not (d244, d164);
	and (d245, d160, d171);
	nor (d246, d164, d204);
	and (d247, d156, d197);
	nand (d248, d158, d176);
	nor (d249, d161, d175);
	nand (d250, d184, d201);
	or (d251, d166, d206);
	nand (d252, d153, d205);
	nor (d253, d175, d206);
	nor (d254, d159, d200);
	buf (d255, d85);
	xnor (d256, d150, d156);
	xor (d257, d184, d207);
	buf (d258, d5);
	and (d259, d157, d186);
	nor (d260, d161, d177);
	nor (d261, d150, d198);
	and (d262, d149, d176);
	nand (d263, d202, d206);
	or (d264, d155, d196);
	or (d265, d152, d187);
	nor (d266, d155, d179);
	buf (d267, d182);
	xor (d268, d176, d190);
	nor (d269, d158, d168);
	xnor (d270, d186, d188);
	and (d271, d154, d168);
	nand (d272, d166, d175);
	xor (d273, d176, d185);
	buf (d274, d110);
	nor (d275, d177, d188);
	nor (d276, d157, d186);
	nor (d277, d162, d170);
	xnor (d278, d162, d189);
	xnor (d279, d172, d187);
	not (d280, d157);
	not (d281, d131);
	not (d282, d110);
	xor (d283, d157, d199);
	nor (d284, d158, d191);
	assign f1 = d280;
	assign f2 = d221;
	assign f3 = d279;
	assign f4 = d241;
endmodule
