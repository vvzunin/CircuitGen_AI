module CCGRCG143( x0, x1, x2, x3, x4, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16 );

	input x0, x1, x2, x3, x4;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290;

	nand (d1, x0, x4);
	nor (d2, x0, x1);
	or (d3, x4);
	xor (d4, x2, x3);
	or (d5, x0);
	not (d6, x2);
	xnor (d7, x2, x3);
	xnor (d8, x2, x4);
	buf (d9, x4);
	xor (d10, x0, x2);
	buf (d11, x1);
	and (d12, x1, x3);
	xor (d13, x3, x4);
	nor (d14, x1, x3);
	xnor (d15, x0, x2);
	and (d16, x4);
	buf (d17, x0);
	and (d18, x1, x3);
	or (d19, x1, x2);
	and (d20, x0, x3);
	and (d21, x0, x3);
	not (d22, x1);
	buf (d23, x2);
	and (d24, x0, x4);
	nor (d25, x0, x4);
	nor (d26, x3, x4);
	xor (d27, x2, x4);
	not (d28, x4);
	xor (d29, x1, x2);
	xor (d30, x0, x1);
	nand (d31, x0);
	nand (d32, x0, x3);
	nand (d33, x3, x4);
	or (d34, x2, x4);
	and (d35, x0, x2);
	nor (d36, x1, x4);
	xor (d37, x2, x3);
	and (d38, x1, x4);
	nand (d39, x1, x4);
	buf (d40, x3);
	xnor (d41, x1, x2);
	not (d42, d1);
	xor (d43, d22, d33);
	and (d44, d11, d39);
	or (d45, d1, d28);
	or (d46, d29, d38);
	xnor (d47, d17, d34);
	xor (d48, d7, d28);
	not (d49, d14);
	and (d50, d19, d40);
	xor (d51, d5, d10);
	xnor (d52, d8, d20);
	buf (d53, d40);
	xnor (d54, d5, d37);
	or (d55, d3, d25);
	xnor (d56, d21, d24);
	xnor (d57, d15, d36);
	not (d58, d22);
	and (d59, d22, d27);
	xor (d60, d11, d22);
	xor (d61, d27, d33);
	xor (d62, d23, d38);
	nand (d63, d14, d19);
	xnor (d64, d14, d23);
	or (d65, d35, d40);
	buf (d66, d22);
	buf (d67, d20);
	nor (d68, d16, d21);
	xnor (d69, d16, d37);
	xor (d70, d29, d40);
	nand (d71, d4, d6);
	nor (d72, d25, d34);
	nor (d73, d29, d32);
	nor (d74, d27, d38);
	and (d75, d13, d24);
	xnor (d76, d5, d15);
	xor (d77, d4, d30);
	and (d78, d4, d25);
	xnor (d79, d11, d35);
	buf (d80, d8);
	or (d81, d11, d23);
	xor (d82, d7, d22);
	buf (d83, d30);
	or (d84, d21, d35);
	xnor (d85, d2, d15);
	buf (d86, d5);
	and (d87, d5, d11);
	xnor (d88, d31, d38);
	and (d89, d11, d33);
	xor (d90, d30, d38);
	or (d91, d12, d15);
	nor (d92, d19, d32);
	not (d93, d15);
	not (d94, d33);
	not (d95, d18);
	buf (d96, d13);
	nor (d97, d5, d12);
	nand (d98, d6, d8);
	xnor (d99, d4, d5);
	nand (d100, d26, d27);
	buf (d101, d19);
	buf (d102, d12);
	or (d103, d4, d11);
	xor (d104, d3, d7);
	nand (d105, d12, d17);
	not (d106, d38);
	or (d107, d16, d20);
	xnor (d108, d11, d26);
	nor (d109, d23, d37);
	not (d110, d40);
	xor (d111, d84, d95);
	nand (d112, d76, d100);
	not (d113, d23);
	and (d114, d61, d83);
	not (d115, d68);
	xor (d116, d96, d100);
	xnor (d117, d60, d65);
	nand (d118, d58, d76);
	nand (d119, d52, d77);
	xnor (d120, d51, d74);
	xnor (d121, d66, d87);
	or (d122, d45, d48);
	xor (d123, d51, d71);
	nor (d124, d75, d95);
	or (d125, d72, d85);
	not (d126, d82);
	nand (d127, d43, d68);
	buf (d128, d81);
	nand (d129, d45, d109);
	buf (d130, d1);
	buf (d131, d21);
	not (d132, d47);
	nor (d133, d63, d70);
	nor (d134, d42, d77);
	buf (d135, d94);
	xor (d136, d62, d109);
	buf (d137, d93);
	nand (d138, d84, d110);
	not (d139, d110);
	nand (d140, d51, d60);
	xor (d141, d57, d97);
	nor (d142, d77, d79);
	and (d143, d96, d102);
	or (d144, d46, d97);
	not (d145, d5);
	or (d146, d88, d108);
	xnor (d147, d54, d64);
	and (d148, d68, d101);
	nor (d149, d73, d80);
	nand (d150, d61, d102);
	nor (d151, d49, d92);
	nor (d152, d67, d82);
	nor (d153, d97, d106);
	not (d154, d67);
	nand (d155, d78, d90);
	and (d156, d45, d109);
	or (d157, d51, d104);
	xor (d158, d46, d60);
	or (d159, d58, d107);
	nor (d160, d69, d91);
	buf (d161, d90);
	or (d162, d48, d87);
	not (d163, d80);
	not (d164, d43);
	xor (d165, d50, d66);
	nor (d166, d63, d104);
	or (d167, d43, d74);
	not (d168, d19);
	or (d169, d76, d84);
	buf (d170, d64);
	buf (d171, d109);
	xnor (d172, d74, d91);
	or (d173, d85, d92);
	not (d174, d86);
	and (d175, d99, d103);
	nand (d176, d48, d55);
	and (d177, d83, d104);
	not (d178, d37);
	or (d179, d142, d165);
	buf (d180, d136);
	xnor (d181, d111, d133);
	nor (d182, d165, d178);
	nand (d183, d150, d169);
	and (d184, d146, d165);
	not (d185, d59);
	or (d186, d164, d168);
	nor (d187, d152, d177);
	nand (d188, d122, d151);
	not (d189, d71);
	and (d190, d137, d152);
	and (d191, d141, d158);
	nor (d192, d130, d177);
	nor (d193, d147, d161);
	and (d194, d116, d163);
	xor (d195, d155, d169);
	and (d196, d116, d117);
	xnor (d197, d143, d161);
	xor (d198, d146, d147);
	and (d199, d133, d143);
	or (d200, d137, d168);
	xnor (d201, d129, d161);
	xor (d202, d164, d173);
	xor (d203, d111, d131);
	nand (d204, d124, d146);
	not (d205, d61);
	not (d206, d96);
	xor (d207, d124, d159);
	xor (d208, d131, d153);
	nor (d209, d162, d169);
	xor (d210, d118, d145);
	xnor (d211, d170, d178);
	xor (d212, d148, d162);
	nor (d213, d111, d112);
	or (d214, d125);
	and (d215, d139, d164);
	nor (d216, d111, d126);
	or (d217, d114, d124);
	xnor (d218, d126, d162);
	and (d219, d132, d163);
	not (d220, d16);
	and (d221, d116, d162);
	xnor (d222, d162, d173);
	not (d223, d12);
	nand (d224, d153, d171);
	nand (d225, d114, d150);
	xor (d226, d142, d168);
	xnor (d227, d129, d174);
	xnor (d228, d123, d165);
	nand (d229, d141, d156);
	not (d230, d128);
	xor (d231, d115, d123);
	nor (d232, d148, d170);
	nor (d233, d141, d155);
	xor (d234, d133, d171);
	buf (d235, d55);
	and (d236, d122, d153);
	xnor (d237, d124, d177);
	and (d238, d143, d158);
	and (d239, d117, d153);
	not (d240, d174);
	xor (d241, d160, d168);
	xnor (d242, d137, d146);
	or (d243, d144, d164);
	not (d244, d84);
	xnor (d245, d137, d139);
	nor (d246, d138, d139);
	nand (d247, d115, d174);
	xnor (d248, d131, d174);
	or (d249, d122, d152);
	not (d250, d8);
	not (d251, d89);
	buf (d252, d63);
	xor (d253, d162, d164);
	nand (d254, d129, d136);
	nand (d255, d135, d159);
	xnor (d256, d153, d166);
	not (d257, d52);
	not (d258, d156);
	and (d259, d118, d133);
	buf (d260, d27);
	and (d261, d117, d138);
	and (d262, d123, d139);
	xor (d263, d147, d149);
	xnor (d264, d122, d136);
	xnor (d265, d197, d201);
	not (d266, d164);
	xor (d267, d225, d235);
	nor (d268, d190, d193);
	and (d269, d181, d200);
	and (d270, d179, d250);
	and (d271, d205, d229);
	nor (d272, d180, d246);
	and (d273, d198, d202);
	nor (d274, d196);
	buf (d275, d135);
	xor (d276, d189, d221);
	nor (d277, d216, d251);
	nor (d278, d191, d194);
	nor (d279, d200, d245);
	nand (d280, d190, d238);
	nand (d281, d199, d200);
	and (d282, d184, d227);
	xor (d283, d210, d252);
	and (d284, d207, d262);
	xor (d285, d222, d253);
	nand (d286, d195, d226);
	buf (d287, d154);
	nand (d288, d240, d245);
	nor (d289, d231, d246);
	nor (d290, d184, d233);
	assign f1 = d272;
	assign f2 = d288;
	assign f3 = d290;
	assign f4 = d272;
	assign f5 = d290;
	assign f6 = d274;
	assign f7 = d286;
	assign f8 = d276;
	assign f9 = d266;
	assign f10 = d279;
	assign f11 = d275;
	assign f12 = d284;
	assign f13 = d268;
	assign f14 = d267;
	assign f15 = d279;
	assign f16 = d290;
endmodule
