module CCGRCG38( x0, x1, x2, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10 );

	input x0, x1, x2;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202;

	or (d1, x0);
	nor (d2, x1, x2);
	not (d3, x1);
	xor (d4, x0, x1);
	buf (d5, x0);
	nor (d6, x2);
	xor (d7, x0, x2);
	nand (d8, x1);
	xor (d9, x1, x2);
	xor (d10, x0);
	or (d11, x0, x2);
	nor (d12, x0);
	and (d13, x0, x2);
	or (d14, x1, x2);
	xor (d15, x1);
	buf (d16, x1);
	and (d17, x2);
	not (d18, x0);
	not (d19, x2);
	xor (d20, x1, x2);
	or (d21, d12, d18);
	buf (d22, d15);
	nand (d23, d10, d12);
	and (d24, d5, d7);
	or (d25, d4, d11);
	buf (d26, d18);
	nand (d27, d5, d17);
	buf (d28, d8);
	buf (d29, d10);
	and (d30, d2, d14);
	nor (d31, d3, d15);
	or (d32, d8, d10);
	not (d33, d8);
	or (d34, d1, d14);
	nor (d35, d18);
	xnor (d36, d1, d4);
	nor (d37, d13, d15);
	and (d38, d6, d17);
	xor (d39, d2, d14);
	not (d40, d3);
	nand (d41, d11, d15);
	not (d42, d14);
	nor (d43, d2, d18);
	or (d44, d4, d12);
	xnor (d45, d12, d18);
	nand (d46, d6, d18);
	and (d47, d1, d15);
	xor (d48, d13, d20);
	or (d49, d6, d14);
	buf (d50, d11);
	xnor (d51, d5, d6);
	buf (d52, d4);
	and (d53, d19, d20);
	nor (d54, d12, d17);
	not (d55, d18);
	xnor (d56, d16, d18);
	or (d57, d11, d12);
	nor (d58, d3, d17);
	xor (d59, d11, d13);
	nand (d60, d21, d39);
	nor (d61, d28, d55);
	and (d62, d33, d34);
	xnor (d63, d26, d49);
	buf (d64, d24);
	and (d65, d48, d50);
	and (d66, d28, d33);
	xor (d67, d60, d66);
	nand (d68, d65);
	xnor (d69, d63, d66);
	nor (d70, d62, d66);
	or (d71, d60, d66);
	or (d72, d63, d64);
	nor (d73, d62);
	and (d74, d61, d62);
	xor (d75, d61, d63);
	not (d76, d55);
	buf (d77, d62);
	or (d78, d62, d63);
	xor (d79, d60, d63);
	buf (d80, d51);
	nand (d81, d62, d65);
	xor (d82, d62, d65);
	nor (d83, d60, d61);
	xor (d84, d63, d66);
	nor (d85, d65, d66);
	and (d86, d62, d63);
	and (d87, d63, d66);
	nand (d88, d63);
	xnor (d89, d60, d64);
	and (d90, d62, d64);
	nand (d91, d62, d66);
	xnor (d92, d61, d64);
	not (d93, d33);
	or (d94, d63, d65);
	and (d95, d62, d63);
	and (d96, d63, d64);
	or (d97, d62, d64);
	not (d98, d57);
	not (d99, d56);
	nand (d100, d60, d62);
	xnor (d101, d60, d61);
	not (d102, d35);
	or (d103, d61, d64);
	not (d104, d32);
	or (d105, d60);
	not (d106, d53);
	nor (d107, d60, d66);
	and (d108, d60, d64);
	xnor (d109, d61, d62);
	buf (d110, d60);
	nor (d111, d64);
	xnor (d112, d63);
	nor (d113, d64, d65);
	not (d114, d36);
	not (d115, d50);
	nor (d116, d65, d66);
	or (d117, d64, d66);
	nand (d118, d64, d65);
	xor (d119, d63, d64);
	nand (d120, d60, d65);
	or (d121, d63);
	xor (d122, d62, d64);
	or (d123, d63, d65);
	nor (d124, d63, d66);
	xor (d125, d60, d61);
	xor (d126, d61, d64);
	xor (d127, d65, d66);
	and (d128, d63);
	buf (d129, d28);
	or (d130, d60, d65);
	xor (d131, d64);
	not (d132, d66);
	xor (d133, d62, d64);
	not (d134, d76);
	and (d135, d71, d84);
	or (d136, d87, d100);
	buf (d137, d91);
	and (d138, d67, d102);
	xor (d139, d104, d111);
	xor (d140, d89, d127);
	nor (d141, d104, d122);
	or (d142, d91, d129);
	xor (d143, d94, d110);
	xor (d144, d84, d126);
	xnor (d145, d136, d140);
	nand (d146, d137, d138);
	xnor (d147, d141, d144);
	xor (d148, d134, d135);
	or (d149, d134, d135);
	xnor (d150, d137);
	nor (d151, d144);
	or (d152, d134, d136);
	buf (d153, d93);
	nor (d154, d139, d140);
	not (d155, d13);
	not (d156, d141);
	or (d157, d139, d144);
	xnor (d158, d135, d142);
	xor (d159, d134, d139);
	xnor (d160, d136, d143);
	xor (d161, d135, d142);
	not (d162, d23);
	not (d163, d2);
	not (d164, d88);
	not (d165, d125);
	nor (d166, d137, d139);
	nor (d167, d135, d138);
	nand (d168, d137, d140);
	xnor (d169, d135);
	or (d170, d143, d144);
	and (d171, d136, d140);
	buf (d172, d2);
	nand (d173, d140);
	nor (d174, d140, d141);
	and (d175, d136, d143);
	nor (d176, d139, d143);
	nand (d177, d135, d142);
	xnor (d178, d136, d142);
	nand (d179, d137, d142);
	nand (d180, d137);
	nor (d181, d134, d138);
	and (d182, d134, d143);
	or (d183, d140, d144);
	xor (d184, d134, d136);
	or (d185, d136, d138);
	xnor (d186, d136, d139);
	or (d187, d143);
	nor (d188, d136, d138);
	nand (d189, d134, d141);
	nand (d190, d135, d136);
	nand (d191, d139, d143);
	xor (d192, d136, d142);
	nor (d193, d136, d140);
	nor (d194, d137, d138);
	xnor (d195, d142, d144);
	and (d196, d142, d143);
	buf (d197, d82);
	nand (d198, d143, d144);
	and (d199, d141, d143);
	and (d200, d138, d141);
	nor (d201, d134, d137);
	and (d202, d134, d144);
	assign f1 = d176;
	assign f2 = d161;
	assign f3 = d148;
	assign f4 = d154;
	assign f5 = d172;
	assign f6 = d186;
	assign f7 = d178;
	assign f8 = d175;
	assign f9 = d197;
	assign f10 = d175;
endmodule
