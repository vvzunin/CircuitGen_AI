module CCGRCG42( x0, x1, x2, f1, f2, f3, f4 );

	input x0, x1, x2;
	output f1, f2, f3, f4;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309;

	xor (d1, x0, x1);
	nand (d2, x1);
	or (d3, x1);
	xor (d4, x1, x2);
	and (d5, x1, x2);
	xnor (d6, x0);
	xor (d7, x0, x1);
	not (d8, x0);
	buf (d9, x2);
	and (d10, x1, x2);
	xor (d11, x1, x2);
	nor (d12, x1);
	or (d13, x0, x2);
	nand (d14, x1, x2);
	nor (d15, x0, x1);
	nor (d16, x0, x2);
	not (d17, x1);
	or (d18, x1, x2);
	and (d19, x0, x2);
	xnor (d20, x0, x2);
	and (d21, x0);
	or (d22, x0, x2);
	or (d23, x2);
	xnor (d24, x1, x2);
	and (d25, x0, x1);
	and (d26, x0, x1);
	xor (d27, x0, x2);
	not (d28, x2);
	xor (d29, x1);
	and (d30, x1);
	xor (d31, x0, x2);
	or (d32, x0, x1);
	xnor (d33, x2);
	buf (d34, x0);
	nand (d35, x1, x2);
	nand (d36, x0, x2);
	xnor (d37, d9, d36);
	or (d38, d8);
	buf (d39, d25);
	xnor (d40, d29, d33);
	xnor (d41, d3, d34);
	or (d42, d1, d18);
	nand (d43, d10, d28);
	nor (d44, d24);
	not (d45, d24);
	and (d46, d5, d24);
	or (d47, d9, d11);
	not (d48, d11);
	not (d49, d1);
	not (d50, d22);
	and (d51, d23, d36);
	nand (d52, d7, d20);
	buf (d53, d31);
	nor (d54, d4);
	nor (d55, d27, d31);
	nor (d56, d13, d15);
	buf (d57, d9);
	nand (d58, d30, d32);
	and (d59, d13, d28);
	xor (d60, d1, d17);
	and (d61, d2, d15);
	and (d62, d9, d30);
	or (d63, d3, d19);
	or (d64, d20, d24);
	nor (d65, d29, d31);
	not (d66, d26);
	nand (d67, d15, d31);
	and (d68, d10, d25);
	or (d69, d22, d23);
	nand (d70, d11, d12);
	and (d71, d29, d34);
	and (d72, d31, d32);
	nor (d73, d10, d25);
	xor (d74, d15, d29);
	xor (d75, d15, d24);
	buf (d76, d15);
	xor (d77, d8, d9);
	buf (d78, d2);
	and (d79, d17, d33);
	xnor (d80, d11, d21);
	xor (d81, d18, d35);
	nand (d82, d15, d34);
	xor (d83, d13, d23);
	and (d84, d28, d35);
	nor (d85, d18, d35);
	xnor (d86, d5, d20);
	nor (d87, d10, d36);
	and (d88, d5, d10);
	xor (d89, d1, d23);
	and (d90, d8, d21);
	nand (d91, d6, d31);
	xor (d92, d14, d21);
	or (d93, d6, d17);
	or (d94, d12, d21);
	xor (d95, d21, d22);
	not (d96, d10);
	and (d97, d23, d33);
	xor (d98, d13, d27);
	xor (d99, d19, d35);
	and (d100, d18, d34);
	not (d101, d51);
	xnor (d102, d54, d85);
	nor (d103, d40, d53);
	buf (d104, d13);
	xnor (d105, d58, d77);
	not (d106, d28);
	xnor (d107, d97, d100);
	buf (d108, d89);
	xor (d109, d60, d61);
	xnor (d110, d97, d98);
	not (d111, d89);
	nor (d112, d71, d93);
	nor (d113, d74, d83);
	nor (d114, d75, d83);
	nand (d115, d49, d89);
	buf (d116, d19);
	buf (d117, d82);
	or (d118, d43, d81);
	not (d119, d48);
	buf (d120, d38);
	and (d121, d46, d80);
	and (d122, d63, d71);
	nand (d123, d53, d67);
	and (d124, d44, d71);
	nor (d125, d50, d92);
	buf (d126, d14);
	not (d127, d70);
	not (d128, d98);
	or (d129, d64, d99);
	xnor (d130, d90, d93);
	nor (d131, d41, d75);
	xor (d132, d40, d53);
	or (d133, d47, d92);
	nor (d134, d38, d85);
	xor (d135, d49, d86);
	xnor (d136, d57, d97);
	xnor (d137, d44, d58);
	not (d138, d99);
	or (d139, d48, d100);
	nand (d140, d43, d91);
	xor (d141, d45, d57);
	and (d142, d50, d88);
	or (d143, d52, d72);
	nand (d144, d71, d87);
	not (d145, d18);
	xnor (d146, d90, d100);
	xor (d147, d62, d78);
	xnor (d148, d43, d71);
	or (d149, d38, d48);
	nor (d150, d46, d100);
	and (d151, d80, d94);
	not (d152, d87);
	nand (d153, d46, d59);
	xnor (d154, d56, d65);
	or (d155, d77, d90);
	buf (d156, d39);
	and (d157, d46, d74);
	or (d158, d55, d93);
	not (d159, d91);
	xnor (d160, d42, d81);
	and (d161, d45, d78);
	xor (d162, d41, d66);
	or (d163, d49);
	and (d164, d46, d88);
	buf (d165, d52);
	nor (d166, d65, d90);
	xnor (d167, d77, d88);
	xnor (d168, d78, d94);
	buf (d169, d6);
	nor (d170, d42, d94);
	and (d171, d70, d78);
	nor (d172, d70, d73);
	and (d173, d51, d73);
	and (d174, d78, d97);
	nand (d175, d47, d48);
	nand (d176, d59, d72);
	nand (d177, d37, d58);
	xnor (d178, d38, d57);
	nor (d179, d58, d82);
	and (d180, d49, d52);
	xnor (d181, d47, d60);
	and (d182, d72, d80);
	nor (d183, d64, d73);
	xor (d184, d41, d76);
	and (d185, d52, d96);
	xnor (d186, d57, d66);
	or (d187, d57, d68);
	xnor (d188, d67, d70);
	or (d189, d50, d88);
	not (d190, d2);
	xor (d191, d63, d83);
	or (d192, d61, d73);
	nor (d193, d55, d68);
	and (d194, d69);
	not (d195, d36);
	xor (d196, d169, d177);
	and (d197, d119, d182);
	or (d198, d119, d151);
	or (d199, d165, d180);
	xor (d200, d117, d190);
	nor (d201, d123, d180);
	buf (d202, d135);
	xnor (d203, d118, d174);
	xor (d204, d103, d107);
	nand (d205, d120, d142);
	nor (d206, d101, d173);
	buf (d207, d188);
	nor (d208, d106, d179);
	nand (d209, d107, d118);
	or (d210, d150, d188);
	nand (d211, d106, d167);
	nand (d212, d155, d164);
	nor (d213, d136, d163);
	or (d214, d124, d143);
	buf (d215, d103);
	not (d216, d155);
	buf (d217, d43);
	and (d218, d103, d122);
	not (d219, d72);
	or (d220, d112, d129);
	and (d221, d119, d157);
	xnor (d222, d115, d179);
	nor (d223, d145, d171);
	and (d224, d148, d153);
	nand (d225, d128, d182);
	nand (d226, d139, d184);
	and (d227, d197, d208);
	xnor (d228, d201, d204);
	nor (d229, d201, d211);
	buf (d230, d209);
	not (d231, d211);
	nor (d232, d224);
	nand (d233, d198, d205);
	nor (d234, d204, d223);
	and (d235, d205, d210);
	xor (d236, d208, d221);
	and (d237, d206, d221);
	xnor (d238, d207, d210);
	xor (d239, d217, d221);
	xnor (d240, d211, d216);
	xor (d241, d208, d223);
	nor (d242, d195, d218);
	and (d243, d207, d211);
	or (d244, d201, d222);
	xnor (d245, d200, d218);
	xnor (d246, d209, d216);
	buf (d247, d60);
	or (d248, d210, d224);
	and (d249, d206, d225);
	nand (d250, d196, d208);
	xor (d251, d218, d222);
	or (d252, d215, d224);
	xnor (d253, d215, d218);
	buf (d254, d176);
	xnor (d255, d196, d212);
	not (d256, d14);
	xnor (d257, d208, d216);
	not (d258, d112);
	xnor (d259, d202, d213);
	or (d260, d207, d215);
	nor (d261, d208, d212);
	xor (d262, d204, d220);
	or (d263, d213, d218);
	and (d264, d199, d200);
	not (d265, d102);
	and (d266, d199, d210);
	buf (d267, d207);
	or (d268, d209, d219);
	or (d269, d201, d203);
	nand (d270, d209, d218);
	xnor (d271, d223, d224);
	not (d272, d107);
	and (d273, d241, d269);
	nand (d274, d231, d248);
	xor (d275, d229, d249);
	xor (d276, d229, d256);
	xnor (d277, d234, d247);
	and (d278, d246, d254);
	buf (d279, d165);
	nor (d280, d247, d261);
	xor (d281, d232, d259);
	nand (d282, d238, d246);
	xnor (d283, d242, d269);
	not (d284, d124);
	buf (d285, d170);
	xor (d286, d249, d262);
	nor (d287, d258, d261);
	xnor (d288, d252, d268);
	and (d289, d257, d271);
	nand (d290, d243, d265);
	or (d291, d230, d234);
	and (d292, d231, d240);
	and (d293, d235, d246);
	nor (d294, d238, d259);
	not (d295, d222);
	nor (d296, d254, d259);
	not (d297, d219);
	nand (d298, d244, d247);
	xnor (d299, d249, d256);
	xnor (d300, d256, d270);
	xnor (d301, d233, d258);
	not (d302, d169);
	or (d303, d237, d242);
	or (d304, d231, d251);
	and (d305, d228, d232);
	xnor (d306, d238, d248);
	nor (d307, d228, d254);
	or (d308, d254, d256);
	buf (d309, d167);
	assign f1 = d272;
	assign f2 = d299;
	assign f3 = d291;
	assign f4 = d273;
endmodule
