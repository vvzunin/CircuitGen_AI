module CCGRCG196( x0, x1, x2, x3, x4, x5, x6, f1, f2, f3, f4, f5 );

	input x0, x1, x2, x3, x4, x5, x6;
	output f1, f2, f3, f4, f5;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314, d315, d316, d317, d318, d319, d320, d321, d322, d323, d324, d325, d326, d327, d328, d329;

	nand (d1, x0, x4);
	and (d2, x2, x3);
	xor (d3, x2);
	nand (d4, x3, x5);
	buf (d5, x6);
	or (d6, x4, x6);
	or (d7, x5, x6);
	xor (d8, x3, x5);
	nor (d9, x0, x4);
	or (d10, x1);
	xor (d11, x1, x2);
	buf (d12, x4);
	xnor (d13, x4, x6);
	buf (d14, x3);
	xnor (d15, x1, x3);
	not (d16, x3);
	xnor (d17, x5);
	nor (d18, x5, x6);
	and (d19, x0, x5);
	xnor (d20, d13, d15);
	xor (d21, d10, d14);
	xor (d22, d2, d7);
	nor (d23, d4, d6);
	not (d24, d15);
	and (d25, d4, d18);
	xor (d26, d5, d7);
	xor (d27, d5, d14);
	buf (d28, d3);
	and (d29, d1, d9);
	xnor (d30, d1, d17);
	and (d31, d5, d18);
	or (d32, d9, d15);
	xnor (d33, d8, d14);
	nand (d34, d10);
	nand (d35, d4, d19);
	or (d36, d10, d16);
	not (d37, d7);
	or (d38, d3, d17);
	not (d39, d19);
	not (d40, d13);
	not (d41, x0);
	nor (d42, d14, d16);
	not (d43, d3);
	buf (d44, x2);
	nand (d45, d7, d14);
	not (d46, x6);
	nand (d47, d9, d11);
	xnor (d48, d8, d11);
	xnor (d49, d46);
	xnor (d50, d27, d43);
	and (d51, d37, d40);
	and (d52, d24, d38);
	xnor (d53, d30, d44);
	xor (d54, d27, d34);
	and (d55, d36, d42);
	and (d56, d24, d40);
	nor (d57, d20, d40);
	buf (d58, d6);
	nand (d59, d22, d31);
	not (d60, d36);
	or (d61, d31, d48);
	or (d62, d32, d39);
	and (d63, d40, d41);
	xor (d64, d25, d34);
	xor (d65, d23, d29);
	xor (d66, d28, d46);
	not (d67, d47);
	nand (d68, d26, d33);
	not (d69, d29);
	xor (d70, d21, d30);
	xor (d71, d22, d34);
	not (d72, d21);
	xnor (d73, d35, d44);
	or (d74, d28, d32);
	or (d75, d43, d45);
	nor (d76, d26, d44);
	and (d77, d43, d44);
	buf (d78, d2);
	xor (d79, d29, d39);
	nor (d80, d32, d36);
	buf (d81, d40);
	nand (d82, d32, d37);
	nor (d83, d30, d36);
	buf (d84, x0);
	xor (d85, d31, d43);
	xnor (d86, d22, d35);
	buf (d87, d45);
	and (d88, d33, d40);
	xnor (d89, d27, d30);
	not (d90, d18);
	nand (d91, d25, d42);
	xnor (d92, d44, d46);
	nor (d93, d26, d31);
	xor (d94, d31, d42);
	nand (d95, d21, d32);
	buf (d96, d17);
	nand (d97, d56, d76);
	and (d98, d75, d92);
	nor (d99, d54, d57);
	not (d100, d6);
	not (d101, d75);
	xor (d102, d68, d78);
	nor (d103, d49, d64);
	or (d104, d55, d63);
	not (d105, d4);
	and (d106, d67, d73);
	not (d107, d61);
	nor (d108, d62, d90);
	and (d109, d66, d77);
	buf (d110, d84);
	xor (d111, d51, d85);
	xnor (d112, d52, d64);
	xnor (d113, d67, d68);
	and (d114, d73, d85);
	or (d115, d54, d58);
	xnor (d116, d63, d89);
	not (d117, d87);
	xnor (d118, d64, d68);
	and (d119, d74, d78);
	and (d120, d64, d91);
	not (d121, d53);
	or (d122, d79, d89);
	xnor (d123, d87, d88);
	xor (d124, d80, d92);
	xnor (d125, d79, d88);
	nor (d126, d51, d81);
	xor (d127, d55, d85);
	not (d128, d42);
	xor (d129, d61, d83);
	xor (d130, d72, d90);
	or (d131, d54, d62);
	and (d132, d54, d95);
	xor (d133, d64, d74);
	or (d134, d58, d77);
	buf (d135, d69);
	buf (d136, x5);
	xor (d137, d58, d81);
	nand (d138, d60, d65);
	or (d139, d59, d78);
	and (d140, d67, d72);
	nand (d141, d63, d73);
	xor (d142, d49, d89);
	buf (d143, d78);
	or (d144, d51, d57);
	buf (d145, d86);
	buf (d146, d54);
	not (d147, d41);
	nor (d148, d64, d77);
	nand (d149, d89, d90);
	xnor (d150, d58, d61);
	nor (d151, d51, d67);
	xor (d152, d80, d95);
	nor (d153, d53, d85);
	xnor (d154, d66, d77);
	buf (d155, d65);
	or (d156, d51, d83);
	nand (d157, d55, d81);
	not (d158, d37);
	nand (d159, d57, d67);
	nand (d160, d74, d88);
	xor (d161, d71, d79);
	and (d162, d69, d80);
	xor (d163, d53, d68);
	and (d164, d65, d85);
	or (d165, d72);
	not (d166, d48);
	buf (d167, d9);
	or (d168, d79, d92);
	or (d169, d67, d87);
	buf (d170, d27);
	nor (d171, d88, d94);
	buf (d172, d12);
	or (d173, d54, d72);
	and (d174, d61, d80);
	nand (d175, d72, d80);
	and (d176, d87, d91);
	xor (d177, d52, d78);
	nor (d178, d138, d159);
	not (d179, d166);
	or (d180, d102, d170);
	xor (d181, d106, d172);
	nor (d182, d145, d161);
	nor (d183, d144, d154);
	and (d184, d182, d183);
	nand (d185, d180, d182);
	not (d186, d131);
	not (d187, d31);
	nor (d188, d186);
	and (d189, d185, d186);
	buf (d190, d164);
	nand (d191, d185);
	and (d192, d184, d186);
	nand (d193, d184, d185);
	buf (d194, d32);
	nor (d195, d185);
	nor (d196, d184, d186);
	xor (d197, d185, d186);
	and (d198, d186);
	xnor (d199, d184, d186);
	buf (d200, d100);
	xnor (d201, d184);
	or (d202, d185, d186);
	buf (d203, d142);
	xnor (d204, d185, d186);
	and (d205, d185, d186);
	nor (d206, d185, d186);
	nand (d207, d184, d185);
	nor (d208, d184, d185);
	buf (d209, d1);
	or (d210, d185);
	xnor (d211, d185, d186);
	nand (d212, d185, d186);
	buf (d213, d117);
	or (d214, d186);
	nand (d215, d184);
	xor (d216, d184, d186);
	or (d217, d184, d185);
	nand (d218, d185, d186);
	xnor (d219, d184, d186);
	xor (d220, d185, d186);
	or (d221, d184, d186);
	nor (d222, d184, d185);
	not (d223, d120);
	nor (d224, d185, d186);
	or (d225, d185, d186);
	nand (d226, d184, d186);
	not (d227, d86);
	buf (d228, d109);
	not (d229, d130);
	buf (d230, d37);
	xor (d231, d184, d185);
	xnor (d232, d184, d185);
	and (d233, d184, d185);
	buf (d234, d140);
	buf (d235, d159);
	not (d236, d54);
	xor (d237, d184, d185);
	not (d238, d59);
	and (d239, d184, d185);
	xor (d240, d185);
	not (d241, d186);
	not (d242, d105);
	buf (d243, d92);
	buf (d244, d14);
	nor (d245, d184, d186);
	xnor (d246, d184, d185);
	not (d247, d14);
	xor (d248, d200, d223);
	not (d249, d146);
	nand (d250, d234, d242);
	and (d251, d192, d195);
	xnor (d252, d211, d238);
	and (d253, d187, d226);
	nand (d254, d194, d200);
	and (d255, d193, d221);
	not (d256, d106);
	nor (d257, d207, d233);
	xor (d258, d210, d244);
	buf (d259, d243);
	buf (d260, d105);
	xor (d261, d187, d216);
	buf (d262, d107);
	not (d263, d119);
	buf (d264, d201);
	nor (d265, d224, d247);
	nor (d266, d187, d238);
	xor (d267, d208, d222);
	nor (d268, d200, d247);
	nand (d269, d212, d229);
	nand (d270, d206, d231);
	xor (d271, d233, d247);
	nand (d272, d187, d212);
	xnor (d273, d237, d242);
	nor (d274, d221, d244);
	nand (d275, d204, d241);
	nand (d276, d210, d220);
	or (d277, d187, d240);
	nor (d278, d188, d193);
	buf (d279, d160);
	and (d280, d200, d210);
	xor (d281, d190, d199);
	buf (d282, d56);
	xnor (d283, d218, d233);
	xnor (d284, d188, d227);
	not (d285, d100);
	and (d286, d219, d239);
	xor (d287, d243, d247);
	nor (d288, d214, d232);
	or (d289, d205, d233);
	xor (d290, d187, d232);
	xor (d291, d193, d208);
	xnor (d292, d230, d241);
	xor (d293, d219, d223);
	and (d294, d191, d229);
	nand (d295, d218, d224);
	not (d296, d188);
	not (d297, d40);
	nor (d298, d225, d239);
	and (d299, d219, d229);
	xor (d300, d221, d231);
	or (d301, d193, d235);
	xnor (d302, d202, d237);
	xor (d303, d194, d233);
	not (d304, d25);
	buf (d305, d212);
	buf (d306, d102);
	buf (d307, d70);
	not (d308, d196);
	nand (d309, d201, d210);
	nand (d310, d214, d234);
	xnor (d311, d214);
	not (d312, d179);
	or (d313, d207, d227);
	buf (d314, d82);
	and (d315, d193, d194);
	nor (d316, d189, d240);
	and (d317, d206, d241);
	xor (d318, d192, d239);
	xor (d319, d222, d230);
	xnor (d320, d204, d217);
	nor (d321, d223, d238);
	buf (d322, d7);
	xor (d323, d214, d235);
	xor (d324, d236, d240);
	xnor (d325, d205, d227);
	nand (d326, d231, d239);
	or (d327, d189, d197);
	xnor (d328, d193, d203);
	and (d329, d212, d242);
	assign f1 = d267;
	assign f2 = d315;
	assign f3 = d309;
	assign f4 = d310;
	assign f5 = d261;
endmodule
