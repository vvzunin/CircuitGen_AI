module CCGRCG25( x0, x1, x2, f1, f2, f3 );

	input x0, x1, x2;
	output f1, f2, f3;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245;

	nand (d1, x0);
	and (d2, x0, x1);
	and (d3, x1, x2);
	nor (d4, x0, x1);
	nand (d5, x1);
	nor (d6, x0, x2);
	not (d7, x1);
	nand (d8, x0, x2);
	buf (d9, x1);
	nor (d10, x1, x2);
	and (d11, x0);
	xor (d12, x0);
	nand (d13, x0, x2);
	xor (d14, x0, x2);
	xor (d15, x2);
	or (d16, x1);
	xor (d17, x1, x2);
	xnor (d18, x0, x1);
	nor (d19, x0, x1);
	xor (d20, x0, x1);
	xnor (d21, x1);
	buf (d22, x0);
	xnor (d23, x0, x2);
	nor (d24, x1, x2);
	not (d25, x0);
	or (d26, x0, x1);
	or (d27, x0);
	or (d28, x0, x2);
	and (d29, x2);
	xnor (d30, x0, x2);
	xor (d31, x1);
	buf (d32, d22);
	and (d33, d18, d21);
	xor (d34, d16, d17);
	buf (d35, d13);
	nand (d36, d14, d23);
	or (d37, d10, d30);
	or (d38, d4, d5);
	and (d39, d5, d12);
	xor (d40, d6, d23);
	nand (d41, d6, d31);
	xor (d42, d8, d28);
	xor (d43, d5, d7);
	or (d44, d4, d26);
	nor (d45, d11, d15);
	or (d46, d25, d31);
	and (d47, d20);
	nor (d48, d12, d24);
	xor (d49, d4, d29);
	and (d50, d19, d25);
	buf (d51, d19);
	nor (d52, d21, d29);
	xor (d53, d6, d12);
	and (d54, d3, d14);
	nor (d55, d13, d17);
	not (d56, d21);
	xnor (d57, d9, d10);
	or (d58, d9, d31);
	nand (d59, d12, d26);
	xnor (d60, d27, d28);
	not (d61, d31);
	xor (d62, d10, d30);
	or (d63, d27);
	nand (d64, d15, d27);
	or (d65, d1, d27);
	xnor (d66, d6, d10);
	nor (d67, d14, d30);
	not (d68, d26);
	xnor (d69, d9, d30);
	not (d70, d4);
	buf (d71, d28);
	or (d72, d17, d29);
	buf (d73, d17);
	nor (d74, d12, d28);
	nor (d75, d10, d18);
	or (d76, d5);
	xnor (d77, d16, d24);
	xor (d78, d7, d23);
	or (d79, d13, d27);
	nor (d80, d26, d29);
	and (d81, d13, d29);
	xor (d82, d2, d9);
	or (d83, d8, d30);
	nor (d84, d21, d31);
	xnor (d85, d15, d23);
	or (d86, d10, d29);
	xor (d87, d8, d12);
	buf (d88, d6);
	xor (d89, d5, d25);
	xor (d90, d6, d15);
	xor (d91, d35, d51);
	nor (d92, d54, d85);
	xnor (d93, d46, d59);
	nand (d94, d58, d82);
	xor (d95, d44, d90);
	buf (d96, d38);
	nor (d97, d37, d84);
	nor (d98, d68, d90);
	nand (d99, d57, d66);
	or (d100, d55, d87);
	xnor (d101, d51, d76);
	xor (d102, d51, d75);
	nor (d103, d52, d80);
	not (d104, d81);
	not (d105, d84);
	nand (d106, d75, d84);
	and (d107, d44, d46);
	nor (d108, d44, d68);
	not (d109, d87);
	nor (d110, d41, d87);
	xor (d111, d66, d88);
	not (d112, d19);
	nand (d113, d58, d61);
	nor (d114, d64, d77);
	not (d115, d82);
	or (d116, d48, d83);
	not (d117, d60);
	nor (d118, d38, d67);
	nand (d119, d33, d63);
	nor (d120, d36, d55);
	nand (d121, d54, d61);
	not (d122, d63);
	xor (d123, d60, d74);
	nand (d124, d47, d49);
	xor (d125, d66, d79);
	and (d126, d62, d64);
	nor (d127, d42, d88);
	not (d128, d6);
	not (d129, d29);
	not (d130, d77);
	xnor (d131, d55, d80);
	not (d132, d54);
	or (d133, d46);
	buf (d134, d74);
	xnor (d135, d46, d70);
	buf (d136, d2);
	and (d137, d55, d88);
	or (d138, d39, d40);
	and (d139, d43, d48);
	not (d140, d45);
	or (d141, d35, d68);
	nand (d142, d41, d79);
	or (d143, d85, d86);
	not (d144, d40);
	xnor (d145, d41, d66);
	not (d146, d28);
	buf (d147, d64);
	xnor (d148, d63, d72);
	xor (d149, d33, d72);
	or (d150, d85, d86);
	nand (d151, d41, d68);
	not (d152, d75);
	or (d153, d42, d82);
	nand (d154, d64, d82);
	and (d155, d65, d84);
	nor (d156, d78, d89);
	or (d157, d59, d81);
	nand (d158, d42, d78);
	or (d159, d65, d85);
	xor (d160, d59, d75);
	and (d161, d49, d57);
	xor (d162, d66, d84);
	not (d163, d1);
	nand (d164, d118, d146);
	xor (d165, d91, d126);
	or (d166, d104, d124);
	xnor (d167, d164);
	or (d168, d163, d166);
	and (d169, d164, d165);
	not (d170, d139);
	not (d171, d85);
	xor (d172, d165);
	not (d173, d97);
	nor (d174, d164, d166);
	nand (d175, d165);
	nand (d176, d164, d165);
	or (d177, d165);
	nand (d178, d165, d166);
	xor (d179, d163, d166);
	nor (d180, d163, d165);
	and (d181, d165, d166);
	nand (d182, d163, d166);
	buf (d183, d87);
	nor (d184, d163, d165);
	and (d185, d164, d166);
	nor (d186, d163);
	or (d187, d165, d166);
	xor (d188, d166);
	xnor (d189, d164, d166);
	nand (d190, d166);
	xor (d191, d164, d165);
	xnor (d192, d163, d165);
	nand (d193, d164, d166);
	and (d194, d163);
	nor (d195, d163, d166);
	nor (d196, d165, d166);
	nand (d197, d164);
	and (d198, d164);
	nand (d199, d163, d164);
	or (d200, d163, d165);
	xor (d201, d165, d166);
	xnor (d202, d164, d165);
	nor (d203, d164, d165);
	not (d204, d138);
	and (d205, d163, d165);
	not (d206, d48);
	xnor (d207, d163, d166);
	nor (d208, d164);
	buf (d209, d34);
	nor (d210, d165);
	and (d211, d164, d165);
	buf (d212, d78);
	or (d213, d164, d166);
	not (d214, d93);
	xnor (d215, d165);
	nor (d216, d166);
	nor (d217, d164, d166);
	buf (d218, d119);
	nor (d219, d163, d166);
	and (d220, d163, d166);
	or (d221, d163);
	buf (d222, d166);
	or (d223, d164, d165);
	and (d224, d163, d165);
	and (d225, d163, d166);
	buf (d226, d50);
	buf (d227, d35);
	xor (d228, d163, d166);
	buf (d229, d164);
	and (d230, d182, d200);
	nor (d231, d189, d214);
	nand (d232, d178, d206);
	and (d233, d186, d225);
	nor (d234, d169, d172);
	xor (d235, d174, d187);
	or (d236, d203, d223);
	xnor (d237, d170, d192);
	xnor (d238, d191, d197);
	buf (d239, d200);
	nand (d240, d218, d229);
	xor (d241, d219);
	xor (d242, d173, d177);
	xnor (d243, d199, d221);
	or (d244, d169, d224);
	buf (d245, d184);
	assign f1 = d237;
	assign f2 = d240;
	assign f3 = d238;
endmodule
