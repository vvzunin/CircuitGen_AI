module CCGRCG159( x0, x1, x2, x3, x4, x5, f1, f2, f3, f4, f5 );

	input x0, x1, x2, x3, x4, x5;
	output f1, f2, f3, f4, f5;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314, d315, d316, d317, d318, d319, d320, d321, d322, d323, d324, d325, d326, d327, d328, d329, d330, d331, d332, d333, d334, d335, d336, d337, d338, d339, d340, d341, d342, d343, d344, d345, d346, d347, d348, d349, d350, d351, d352, d353, d354, d355, d356, d357, d358, d359, d360, d361, d362, d363, d364, d365, d366, d367, d368, d369, d370, d371, d372, d373, d374, d375, d376, d377, d378, d379, d380, d381, d382, d383, d384, d385, d386, d387, d388, d389, d390, d391, d392, d393, d394, d395, d396, d397, d398, d399, d400, d401, d402, d403, d404, d405, d406, d407, d408, d409, d410, d411, d412, d413, d414, d415, d416, d417, d418, d419, d420, d421, d422, d423, d424, d425, d426, d427, d428, d429, d430, d431, d432, d433;

	xnor (d1, x2, x4);
	buf (d2, x5);
	nand (d3, x2, x3);
	not (d4, x5);
	not (d5, x2);
	buf (d6, x1);
	xnor (d7, x3, x4);
	not (d8, x3);
	xnor (d9, x0, x4);
	not (d10, x4);
	and (d11, x1, x2);
	xor (d12, x0);
	xnor (d13, x2);
	and (d14, x3);
	or (d15, x3, x5);
	xnor (d16, x1, x3);
	buf (d17, x2);
	and (d18, x1, x4);
	nand (d19, x0);
	xnor (d20, x1, x4);
	and (d21, x2, x5);
	nand (d22, x0, x3);
	xor (d23, x2, x5);
	xor (d24, x0, x4);
	nor (d25, x0, x3);
	xor (d26, x3, x4);
	nand (d27, x0, x1);
	xnor (d28, x0, x5);
	nor (d29, x1, x4);
	not (d30, x0);
	xor (d31, x1, x4);
	xor (d32, x0, x1);
	nor (d33, x3);
	nand (d34, x2, x4);
	and (d35, x1, x5);
	nor (d36, x0, x2);
	xnor (d37, x2, x3);
	not (d38, x1);
	buf (d39, d23);
	not (d40, d2);
	not (d41, d29);
	nand (d42, d11, d32);
	xnor (d43, d11, d37);
	xor (d44, d23, d38);
	and (d45, d32, d38);
	xnor (d46, d18, d28);
	nand (d47, d32, d36);
	and (d48, d4, d38);
	xor (d49, d3, d32);
	nand (d50, d20, d23);
	buf (d51, d27);
	xor (d52, d2, d4);
	xnor (d53, d5, d27);
	xnor (d54, d4, d23);
	xor (d55, d14, d37);
	nor (d56, d13, d25);
	or (d57, d5, d25);
	or (d58, d8, d19);
	and (d59, d20, d32);
	not (d60, d6);
	not (d61, d22);
	xor (d62, d14, d19);
	xnor (d63, d27, d38);
	nor (d64, d27, d28);
	xnor (d65, d12);
	nor (d66, d21, d33);
	or (d67, d11, d28);
	nand (d68, d36, d38);
	and (d69, d18, d30);
	nor (d70, d7);
	not (d71, d3);
	buf (d72, d13);
	nand (d73, d5, d34);
	nand (d74, d23, d28);
	nand (d75, d25, d30);
	nor (d76, d13, d34);
	or (d77, d7, d14);
	nor (d78, d10, d22);
	nand (d79, d23, d36);
	buf (d80, d36);
	xor (d81, d26, d28);
	nor (d82, d26, d36);
	and (d83, d14, d20);
	not (d84, d19);
	nor (d85, d3, d19);
	nor (d86, d5, d8);
	xor (d87, d4, d34);
	xor (d88, d3, d9);
	or (d89, d58, d69);
	xor (d90, d39, d84);
	and (d91, d48, d49);
	nand (d92, d49, d55);
	nand (d93, d65, d67);
	or (d94, d45, d74);
	xor (d95, d46, d78);
	and (d96, d53, d73);
	nor (d97, d55, d85);
	and (d98, d39, d40);
	buf (d99, d76);
	buf (d100, d50);
	not (d101, d15);
	or (d102, d39, d47);
	nand (d103, d41, d64);
	nand (d104, d64, d77);
	nand (d105, d58, d70);
	xnor (d106, d66, d85);
	not (d107, d51);
	or (d108, d44, d53);
	buf (d109, d69);
	nor (d110, d46, d77);
	buf (d111, d57);
	not (d112, d55);
	nor (d113, d47, d74);
	nand (d114, d63, d79);
	nor (d115, d44, d56);
	xnor (d116, d39, d53);
	and (d117, d60, d74);
	xnor (d118, d56, d61);
	xor (d119, d54, d83);
	nor (d120, d51, d82);
	not (d121, d18);
	nor (d122, d72, d79);
	xnor (d123, d46, d72);
	or (d124, d76, d79);
	and (d125, d42, d59);
	nand (d126, d55, d88);
	xnor (d127, d57, d84);
	xnor (d128, d54, d67);
	not (d129, d33);
	nand (d130, d43, d61);
	nand (d131, d42, d76);
	xor (d132, d40, d88);
	xnor (d133, d41, d73);
	xor (d134, d43, d54);
	buf (d135, d75);
	xnor (d136, d48, d60);
	nor (d137, d55, d81);
	or (d138, d47, d77);
	nor (d139, d52, d80);
	xnor (d140, d43, d74);
	or (d141, d53, d66);
	xor (d142, d59, d84);
	and (d143, d50, d54);
	nand (d144, d53, d67);
	xor (d145, d64, d81);
	nor (d146, d67, d88);
	nor (d147, d57, d69);
	or (d148, d79, d87);
	nor (d149, d57, d75);
	buf (d150, d28);
	xor (d151, d43, d70);
	xnor (d152, d72, d80);
	buf (d153, d55);
	not (d154, d52);
	xor (d155, d70, d80);
	not (d156, d8);
	xnor (d157, d50, d80);
	not (d158, d23);
	buf (d159, d45);
	and (d160, d95, d107);
	xnor (d161, d92, d130);
	buf (d162, d89);
	nor (d163, d113, d117);
	not (d164, d152);
	xnor (d165, d110, d150);
	xnor (d166, d118, d125);
	xor (d167, d122, d127);
	nor (d168, d121, d152);
	xnor (d169, d119, d121);
	or (d170, d106, d115);
	xor (d171, d110, d113);
	and (d172, d143, d149);
	nand (d173, d111, d116);
	nor (d174, d99, d156);
	nor (d175, d97, d108);
	xor (d176, d124, d142);
	xor (d177, d97, d116);
	nand (d178, d119, d129);
	nor (d179, d133, d135);
	xnor (d180, d104, d112);
	xor (d181, d137, d142);
	nor (d182, d99, d119);
	nor (d183, d125, d135);
	xor (d184, d102, d153);
	nand (d185, d145, d152);
	xor (d186, d131, d132);
	xor (d187, d109, d113);
	xnor (d188, d129, d134);
	nor (d189, d128, d135);
	xnor (d190, d91, d139);
	xor (d191, d93, d136);
	or (d192, d107, d146);
	xor (d193, d89, d133);
	and (d194, d122, d144);
	nor (d195, d101, d121);
	nand (d196, d119, d142);
	or (d197, d108, d116);
	nor (d198, d105, d144);
	nor (d199, d91, d124);
	and (d200, d100, d113);
	not (d201, d49);
	nor (d202, d92, d95);
	and (d203, d93, d157);
	and (d204, d129, d136);
	nor (d205, d95, d143);
	nand (d206, d97, d140);
	not (d207, d136);
	not (d208, d92);
	and (d209, d133, d150);
	not (d210, d149);
	xor (d211, d106, d157);
	and (d212, d138, d155);
	nor (d213, d107, d119);
	xor (d214, d125, d153);
	nor (d215, d179, d197);
	not (d216, d209);
	xnor (d217, d199, d209);
	nor (d218, d208, d211);
	xnor (d219, d205, d209);
	and (d220, d180, d189);
	nor (d221, d183, d184);
	or (d222, d165, d181);
	xnor (d223, d191, d208);
	nand (d224, d169, d184);
	and (d225, d165, d198);
	xnor (d226, d160, d206);
	xnor (d227, d193, d210);
	xor (d228, d176, d194);
	not (d229, d153);
	xor (d230, d178, d180);
	not (d231, d167);
	and (d232, d179, d186);
	xnor (d233, d179, d193);
	nor (d234, d175, d185);
	nand (d235, d206, d211);
	buf (d236, d154);
	nor (d237, d172, d179);
	and (d238, d165, d180);
	xnor (d239, d192, d206);
	nor (d240, d191, d203);
	nand (d241, d177, d212);
	not (d242, d46);
	or (d243, d183, d206);
	nor (d244, d187, d204);
	or (d245, d188, d194);
	xnor (d246, d188, d190);
	xnor (d247, d196, d205);
	buf (d248, d48);
	not (d249, d112);
	nor (d250, d172, d202);
	xnor (d251, d164, d201);
	nor (d252, d176, d198);
	nand (d253, d203, d212);
	nor (d254, d185, d198);
	and (d255, d163, d185);
	nor (d256, d198, d213);
	or (d257, d183, d196);
	xor (d258, d172, d178);
	or (d259, d159, d197);
	nand (d260, d173, d187);
	buf (d261, d87);
	xor (d262, d190, d207);
	nand (d263, d163, d199);
	or (d264, d167, d176);
	nor (d265, d171, d195);
	nor (d266, d182, d199);
	or (d267, d173, d189);
	not (d268, d176);
	buf (d269, d184);
	nor (d270, d170, d180);
	xnor (d271, d184, d196);
	nand (d272, d206, d214);
	or (d273, d161, d182);
	nor (d274, d174, d194);
	and (d275, d164, d196);
	and (d276, d159, d206);
	not (d277, d31);
	xnor (d278, d170, d201);
	xnor (d279, d179, d213);
	or (d280, d184, d209);
	xor (d281, d183, d194);
	xnor (d282, d180, d198);
	or (d283, d159, d192);
	and (d284, d163, d174);
	or (d285, d161, d176);
	xor (d286, d169, d188);
	not (d287, d17);
	nand (d288, d193, d211);
	nand (d289, d232, d234);
	xnor (d290, d234, d288);
	xnor (d291, d287);
	xor (d292, d248, d253);
	xnor (d293, d266, d270);
	xor (d294, d243, d276);
	or (d295, d246, d280);
	nand (d296, d232, d254);
	buf (d297, d78);
	xnor (d298, d255, d261);
	xnor (d299, d215, d270);
	buf (d300, d266);
	xnor (d301, d242, d270);
	xnor (d302, d244, d252);
	xnor (d303, d276, d284);
	xor (d304, d220, d237);
	not (d305, d254);
	nand (d306, d238, d266);
	and (d307, d245, d255);
	and (d308, d215, d255);
	nor (d309, d215);
	and (d310, d242, d284);
	xnor (d311, d233, d270);
	and (d312, d221, d247);
	not (d313, d166);
	or (d314, d225, d249);
	xnor (d315, d218, d230);
	or (d316, d256, d257);
	nand (d317, d229, d250);
	buf (d318, d201);
	nor (d319, d220, d261);
	xnor (d320, d234, d284);
	and (d321, d259, d286);
	nand (d322, d233, d248);
	xnor (d323, d244, d277);
	nor (d324, d246, d264);
	and (d325, d249, d281);
	xnor (d326, d225, d257);
	nand (d327, d238, d285);
	buf (d328, d244);
	and (d329, d224, d267);
	xnor (d330, d250, d286);
	xor (d331, d263, d286);
	not (d332, d109);
	nor (d333, d232, d262);
	and (d334, d248, d288);
	or (d335, d244, d259);
	xnor (d336, d219, d286);
	nor (d337, d239, d253);
	or (d338, d222, d243);
	nor (d339, d232, d284);
	not (d340, d86);
	buf (d341, d191);
	xor (d342, d254, d265);
	not (d343, d205);
	not (d344, d264);
	nor (d345, d247, d285);
	xnor (d346, d245, d264);
	nor (d347, d245, d269);
	and (d348, d273, d275);
	xnor (d349, d241, d244);
	buf (d350, d47);
	or (d351, d276, d281);
	nor (d352, d221, d236);
	not (d353, d160);
	or (d354, d217, d282);
	buf (d355, d96);
	not (d356, d227);
	xor (d357, d257, d281);
	or (d358, d248, d258);
	nand (d359, d236, d286);
	and (d360, d250, d281);
	and (d361, d243, d256);
	buf (d362, d282);
	xor (d363, d266, d285);
	not (d364, d131);
	and (d365, d269, d279);
	nand (d366, d235, d240);
	xor (d367, d219, d222);
	nor (d368, d266, d280);
	or (d369, d230, d238);
	and (d370, d244, d261);
	nand (d371, d219, d264);
	xor (d372, d226, d268);
	nor (d373, d238, d275);
	xnor (d374, d245, d248);
	or (d375, d246, d272);
	nor (d376, d221, d263);
	xnor (d377, d226, d251);
	nand (d378, d230, d285);
	not (d379, d162);
	xor (d380, d245, d274);
	xnor (d381, d367, d368);
	not (d382, d317);
	xor (d383, d339, d343);
	nor (d384, d292, d369);
	xnor (d385, d332, d333);
	xor (d386, d341, d353);
	buf (d387, d314);
	nand (d388, d329, d367);
	nand (d389, d331, d379);
	xnor (d390, d383, d389);
	and (d391, d384, d387);
	nand (d392, d388);
	and (d393, d381, d384);
	nor (d394, d381, d384);
	and (d395, d382, d389);
	nor (d396, d385, d389);
	or (d397, d382, d388);
	buf (d398, d149);
	nand (d399, d384, d389);
	xnor (d400, d385, d389);
	nand (d401, d381, d382);
	nand (d402, d384, d385);
	buf (d403, d152);
	buf (d404, d275);
	not (d405, d368);
	buf (d406, d210);
	and (d407, d381, d386);
	buf (d408, d52);
	not (d409, d27);
	xor (d410, d382, d386);
	xor (d411, d383, d385);
	not (d412, d14);
	nor (d413, d385, d387);
	and (d414, d385, d387);
	not (d415, d305);
	nand (d416, d386, d388);
	buf (d417, d254);
	not (d418, d164);
	nand (d419, d382, d383);
	not (d420, d95);
	nand (d421, d385, d388);
	nor (d422, d386, d389);
	nor (d423, d382, d388);
	xor (d424, d383, d385);
	nor (d425, d383, d389);
	xor (d426, d382, d389);
	xnor (d427, d385, d387);
	or (d428, d386, d387);
	and (d429, d382, d385);
	nand (d430, d387, d389);
	xor (d431, d388, d389);
	or (d432, d382, d384);
	xor (d433, d382, d387);
	assign f1 = d392;
	assign f2 = d420;
	assign f3 = d428;
	assign f4 = d422;
	assign f5 = d413;
endmodule
