module CCGRCG150( x0, x1, x2, x3, x4, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17, f18, f19, f20 );

	input x0, x1, x2, x3, x4;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17, f18, f19, f20;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291;

	nand (d1, x0);
	xnor (d2, x3);
	xor (d3, x0, x1);
	xor (d4, x1, x4);
	xnor (d5, x1, x4);
	nor (d6, x3, x4);
	xor (d7, x0, x2);
	or (d8, x3, x4);
	or (d9, x0, x4);
	or (d10, x2, x3);
	xnor (d11, x0, x4);
	or (d12, x2, x4);
	nor (d13, x1);
	buf (d14, x1);
	and (d15, x0, x2);
	buf (d16, x2);
	not (d17, x2);
	and (d18, x3, x4);
	nand (d19, x2);
	buf (d20, x0);
	and (d21, x0, x4);
	or (d22, x0, x2);
	or (d23, x0, x1);
	or (d24, x2, x4);
	not (d25, x3);
	buf (d26, x4);
	and (d27, x0, x4);
	xnor (d28, x0, x1);
	nand (d29, x0, x2);
	xor (d30, x3, x4);
	or (d31, x1, x4);
	xor (d32, x0, x1);
	xor (d33, x1, x3);
	xor (d34, x2, x3);
	buf (d35, x3);
	nand (d36, x2, x4);
	and (d37, x3);
	xnor (d38, x4);
	and (d39, x0, x1);
	xnor (d40, x2, x3);
	nor (d41, x1, x2);
	nand (d42, x0, x1);
	and (d43, x1, x3);
	not (d44, x4);
	not (d45, x0);
	and (d46, x0, x2);
	or (d47, x4);
	nor (d48, x2, x3);
	nand (d49, x0, x4);
	nor (d50, x3);
	nor (d51, x1, x3);
	xor (d52, x0, x4);
	and (d53, d25, d37);
	or (d54, d14, d48);
	xnor (d55, d33, d37);
	nand (d56, d19, d34);
	buf (d57, d28);
	nor (d58, d6, d16);
	and (d59, d4, d34);
	or (d60, d12, d50);
	xor (d61, d12, d43);
	nand (d62, d44, d46);
	xor (d63, d22, d32);
	or (d64, d13, d23);
	nand (d65, d38, d41);
	nor (d66, d19, d32);
	nand (d67, d19, d36);
	xor (d68, d15, d26);
	xnor (d69, d33, d37);
	buf (d70, d45);
	and (d71, d26, d42);
	xnor (d72, d43, d46);
	not (d73, d36);
	buf (d74, d43);
	nor (d75, d29, d35);
	buf (d76, d51);
	or (d77, d42, d43);
	xnor (d78, d38, d50);
	or (d79, d15, d36);
	and (d80, d1, d2);
	or (d81, d27, d48);
	nand (d82, d13, d23);
	nand (d83, d5, d44);
	not (d84, d31);
	and (d85, d43, d48);
	xor (d86, d32, d37);
	not (d87, d46);
	nor (d88, d28, d37);
	not (d89, d18);
	xnor (d90, d19);
	or (d91, d6, d29);
	xnor (d92, d28, d52);
	nand (d93, d5, d43);
	not (d94, d10);
	xor (d95, d13, d31);
	buf (d96, d11);
	nand (d97, d22, d29);
	nor (d98, d1, d37);
	buf (d99, d29);
	xnor (d100, d23, d42);
	buf (d101, d18);
	or (d102, d3, d17);
	xnor (d103, d1, d43);
	buf (d104, d31);
	nand (d105, d17, d31);
	buf (d106, d40);
	nand (d107, d10, d41);
	or (d108, d11, d41);
	not (d109, d27);
	and (d110, d11, d37);
	xnor (d111, d12, d22);
	and (d112, d35, d44);
	nand (d113, d17, d33);
	or (d114, d20, d40);
	buf (d115, d37);
	nand (d116, d4, d12);
	nand (d117, d13, d44);
	nand (d118, d12, d25);
	xnor (d119, d24, d34);
	and (d120, d19, d51);
	not (d121, d51);
	nor (d122, d4, d30);
	not (d123, d49);
	nand (d124, d35, d50);
	xor (d125, d5, d44);
	xnor (d126, d12, d40);
	nor (d127, d4, d18);
	buf (d128, d5);
	and (d129, d2, d39);
	not (d130, d37);
	nor (d131, d103, d123);
	not (d132, d58);
	and (d133, d77, d104);
	xnor (d134, d79, d105);
	buf (d135, d60);
	nand (d136, d60, d126);
	and (d137, d59, d67);
	xnor (d138, d57, d59);
	xor (d139, d84, d90);
	nor (d140, d60, d116);
	xnor (d141, d60, d85);
	nand (d142, d74, d126);
	xor (d143, d55, d109);
	nor (d144, d60, d80);
	and (d145, d90, d124);
	xor (d146, d100, d110);
	nor (d147, d66, d123);
	and (d148, d67, d128);
	nor (d149, d72, d124);
	or (d150, d101, d107);
	xnor (d151, d75, d78);
	not (d152, d24);
	nor (d153, d119, d126);
	not (d154, d80);
	not (d155, d15);
	or (d156, d66, d68);
	buf (d157, d26);
	or (d158, d85, d104);
	buf (d159, d65);
	nor (d160, d53, d127);
	nor (d161, d62, d69);
	not (d162, d100);
	xor (d163, d75, d114);
	xnor (d164, d93, d96);
	xor (d165, d124, d129);
	xor (d166, d82, d105);
	not (d167, d126);
	nand (d168, d55, d98);
	xor (d169, d61, d107);
	xor (d170, d63, d119);
	xor (d171, d69, d113);
	and (d172, d79, d129);
	buf (d173, d63);
	buf (d174, d79);
	or (d175, d161, d166);
	nor (d176, d138, d145);
	and (d177, d135, d155);
	buf (d178, d70);
	xnor (d179, d138, d170);
	or (d180, d140, d161);
	and (d181, d144, d150);
	buf (d182, d170);
	xnor (d183, d143, d168);
	nor (d184, d163, d170);
	or (d185, d142, d168);
	xor (d186, d138, d164);
	buf (d187, d25);
	nor (d188, d132, d152);
	not (d189, d97);
	and (d190, d174, d179);
	nand (d191, d175, d189);
	and (d192, d184, d189);
	xnor (d193, d177, d187);
	and (d194, d175, d180);
	nand (d195, d180, d185);
	nor (d196, d178, d185);
	and (d197, d178, d180);
	nor (d198, d179, d182);
	and (d199, d180);
	nor (d200, d174, d186);
	and (d201, d179);
	and (d202, d178, d185);
	xor (d203, d174, d180);
	nor (d204, d173, d180);
	nor (d205, d178, d179);
	xor (d206, d176, d177);
	and (d207, d173, d188);
	buf (d208, d24);
	xor (d209, d180, d184);
	xnor (d210, d174, d189);
	buf (d211, d17);
	nand (d212, d176, d185);
	nor (d213, d183, d187);
	nor (d214, d180, d182);
	xor (d215, d178, d187);
	nor (d216, d180, d183);
	and (d217, d175, d181);
	and (d218, d185, d187);
	not (d219, d135);
	nand (d220, d174, d180);
	xnor (d221, d173, d174);
	and (d222, d177, d183);
	or (d223, d178, d187);
	nor (d224, d184);
	not (d225, d41);
	buf (d226, d103);
	nand (d227, d178, d185);
	nor (d228, d181, d187);
	xnor (d229, d174, d182);
	not (d230, d121);
	nor (d231, d187, d188);
	xor (d232, d176, d180);
	xnor (d233, d179, d184);
	xnor (d234, d176, d185);
	nor (d235, d179, d186);
	not (d236, d94);
	buf (d237, d148);
	buf (d238, d56);
	buf (d239, d104);
	buf (d240, d121);
	buf (d241, d3);
	xnor (d242, d177, d188);
	nor (d243, d173, d177);
	buf (d244, d82);
	not (d245, d81);
	buf (d246, d157);
	nor (d247, d178, d183);
	not (d248, d3);
	or (d249, d175, d186);
	or (d250, d183, d185);
	xnor (d251, d184, d185);
	and (d252, d178, d188);
	buf (d253, d107);
	nor (d254, d175, d177);
	buf (d255, d146);
	xnor (d256, d176, d179);
	or (d257, d185, d186);
	xnor (d258, d223, d241);
	nor (d259, d193, d247);
	not (d260, d144);
	nand (d261, d193, d195);
	and (d262, d229, d240);
	xor (d263, d246, d257);
	nand (d264, d204, d218);
	xor (d265, d228, d231);
	nand (d266, d209, d243);
	and (d267, d195, d237);
	not (d268, d197);
	or (d269, d238, d252);
	not (d270, d40);
	xor (d271, d209, d234);
	and (d272, d206, d236);
	or (d273, d202, d233);
	xnor (d274, d208, d241);
	xor (d275, d208, d236);
	nor (d276, d209, d252);
	buf (d277, d253);
	buf (d278, d113);
	buf (d279, d187);
	nand (d280, d234, d246);
	xor (d281, d194, d246);
	buf (d282, d13);
	xor (d283, d206, d237);
	xor (d284, d236);
	not (d285, d137);
	xor (d286, d194, d224);
	and (d287, d216, d244);
	not (d288, d63);
	not (d289, d85);
	and (d290, d249, d252);
	xnor (d291, d228, d257);
	assign f1 = d263;
	assign f2 = d291;
	assign f3 = d274;
	assign f4 = d265;
	assign f5 = d265;
	assign f6 = d258;
	assign f7 = d268;
	assign f8 = d261;
	assign f9 = d281;
	assign f10 = d287;
	assign f11 = d263;
	assign f12 = d263;
	assign f13 = d281;
	assign f14 = d279;
	assign f15 = d278;
	assign f16 = d279;
	assign f17 = d278;
	assign f18 = d274;
	assign f19 = d273;
	assign f20 = d281;
endmodule
