module CCGRCG7( x0, x1, f1, f2, f3, f4 );

	input x0, x1;
	output f1, f2, f3, f4;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314, d315, d316, d317, d318, d319, d320, d321, d322, d323, d324, d325, d326, d327, d328, d329, d330, d331, d332, d333, d334, d335, d336, d337, d338, d339, d340, d341, d342, d343, d344, d345, d346, d347, d348, d349, d350, d351, d352, d353, d354, d355, d356;

	xor (d1, x0, x1);
	xor (d2, x0, x1);
	nor (d3, x0, x1);
	and (d4, x0, x1);
	not (d5, x0);
	not (d6, x1);
	buf (d7, x1);
	or (d8, x0, x1);
	nor (d9, x0);
	xnor (d10, x0, x1);
	and (d11, x0, x1);
	or (d12, x0, x1);
	xnor (d13, x0, x1);
	or (d14, x1);
	or (d15, x0);
	nand (d16, x0, x1);
	buf (d17, x0);
	nand (d18, x0, x1);
	nand (d19, x1);
	nor (d20, x0, x1);
	nand (d21, x0);
	xnor (d22, x1);
	and (d23, x0);
	xor (d24, x0);
	nand (d25, d1, d19);
	xnor (d26, d8, d10);
	or (d27, d13, d20);
	not (d28, d9);
	nor (d29, d14, d21);
	or (d30, d12, d15);
	nand (d31, d15, d22);
	buf (d32, d17);
	nor (d33, d16, d17);
	nand (d34, d1, d18);
	or (d35, d6, d14);
	or (d36, d10, d12);
	buf (d37, d19);
	nor (d38, d12, d14);
	and (d39, d2, d16);
	xnor (d40, d2, d6);
	xor (d41, d20, d21);
	nor (d42, d1, d22);
	not (d43, d21);
	xnor (d44, d12, d21);
	xnor (d45, d6, d22);
	xor (d46, d7, d21);
	nor (d47, d11, d23);
	buf (d48, d15);
	nor (d49, d8, d22);
	xor (d50, d10, d13);
	xor (d51, d5, d14);
	and (d52, d3, d22);
	xnor (d53, d13, d22);
	nand (d54, d2, d20);
	and (d55, d14, d16);
	xor (d56, d4, d5);
	xor (d57, d3, d20);
	or (d58, d4, d10);
	or (d59, d10, d12);
	xnor (d60, d10, d16);
	xnor (d61, d3, d14);
	xor (d62, d6, d11);
	nor (d63, d2, d6);
	not (d64, d7);
	and (d65, d13);
	and (d66, d5, d14);
	xnor (d67, d9, d11);
	nand (d68, d12);
	xnor (d69, d6, d16);
	buf (d70, d8);
	or (d71, d10, d14);
	or (d72, d1, d23);
	buf (d73, d24);
	not (d74, d2);
	nand (d75, d20);
	nor (d76, d5, d6);
	xor (d77, d19, d21);
	xor (d78, d1, d12);
	and (d79, d4, d19);
	xor (d80, d12, d19);
	and (d81, d12, d20);
	or (d82, d15, d18);
	and (d83, d5, d7);
	not (d84, d1);
	xnor (d85, d4, d15);
	buf (d86, d10);
	nand (d87, d6, d22);
	xnor (d88, d10, d13);
	nor (d89, d15, d20);
	not (d90, d14);
	and (d91, d3, d6);
	and (d92, d1, d24);
	not (d93, d18);
	xor (d94, d10, d14);
	xnor (d95, d16, d21);
	and (d96, d5, d21);
	and (d97, d8, d11);
	nand (d98, d8, d16);
	and (d99, d12, d23);
	and (d100, d15, d23);
	not (d101, d8);
	nand (d102, d9, d23);
	not (d103, d69);
	nor (d104, d73, d89);
	not (d105, d97);
	not (d106, d74);
	or (d107, d25, d92);
	and (d108, d33, d82);
	xnor (d109, d27, d82);
	nand (d110, d51, d79);
	nand (d111, d62, d66);
	nor (d112, d32, d63);
	or (d113, d78, d94);
	xnor (d114, d29, d83);
	nor (d115, d28, d74);
	and (d116, d37, d54);
	nor (d117, d25, d51);
	or (d118, d105, d109);
	not (d119, d87);
	nor (d120, d112);
	not (d121, d68);
	buf (d122, d65);
	not (d123, d27);
	nand (d124, d114);
	nand (d125, d103, d116);
	or (d126, d116, d117);
	xnor (d127, d111, d116);
	xnor (d128, d113, d114);
	nor (d129, d105, d106);
	buf (d130, d104);
	and (d131, d104, d111);
	nor (d132, d109, d110);
	and (d133, d113, d115);
	nor (d134, d108, d111);
	or (d135, d107, d113);
	not (d136, d43);
	and (d137, d106, d107);
	nor (d138, d107, d114);
	xor (d139, d115);
	not (d140, d28);
	nor (d141, d105, d108);
	nor (d142, d112, d115);
	xor (d143, d103, d117);
	or (d144, d106, d111);
	xor (d145, d114, d115);
	nand (d146, d115);
	buf (d147, d62);
	and (d148, d107, d109);
	xor (d149, d108, d113);
	nand (d150, d106, d107);
	and (d151, d105, d108);
	nor (d152, d103, d109);
	or (d153, d106, d107);
	xor (d154, d106, d108);
	nor (d155, d104, d112);
	and (d156, d108, d111);
	not (d157, d66);
	nor (d158, d104, d117);
	and (d159, d107, d111);
	xor (d160, d103, d106);
	nand (d161, d103, d110);
	buf (d162, d71);
	buf (d163, d103);
	not (d164, d65);
	nand (d165, d106, d114);
	nand (d166, d110, d117);
	and (d167, d105, d106);
	xnor (d168, d108, d117);
	or (d169, d107, d115);
	buf (d170, d25);
	xor (d171, d107, d111);
	xnor (d172, d113, d117);
	nand (d173, d105, d114);
	or (d174, d111, d112);
	not (d175, d78);
	and (d176, d111, d115);
	nor (d177, d112, d116);
	buf (d178, d61);
	or (d179, d107, d116);
	nand (d180, d178, d179);
	or (d181, d136, d161);
	xnor (d182, d140, d175);
	buf (d183, d33);
	and (d184, d119, d146);
	or (d185, d176, d179);
	not (d186, d62);
	not (d187, d164);
	nor (d188, d158, d171);
	and (d189, d151, d166);
	xnor (d190, d121, d130);
	xnor (d191, d118, d158);
	xnor (d192, d125, d145);
	xor (d193, d124, d176);
	xnor (d194, d142, d161);
	xnor (d195, d130, d177);
	not (d196, d116);
	nand (d197, d157, d164);
	nor (d198, d135, d141);
	nor (d199, d120, d137);
	xnor (d200, d160, d168);
	xnor (d201, d153, d161);
	xnor (d202, d130, d157);
	and (d203, d120, d170);
	and (d204, d147, d169);
	xnor (d205, d170);
	xor (d206, d124, d144);
	nor (d207, d118, d133);
	nand (d208, d137, d172);
	xnor (d209, d162, d178);
	xnor (d210, d129, d155);
	nor (d211, d167, d168);
	nand (d212, d122, d137);
	nor (d213, d120, d128);
	buf (d214, d79);
	not (d215, d170);
	xnor (d216, d156, d176);
	nand (d217, d153, d166);
	nand (d218, d129, d168);
	xnor (d219, d141, d148);
	xnor (d220, d155, d164);
	xnor (d221, d118, d139);
	nor (d222, d140, d159);
	nand (d223, d119, d147);
	or (d224, d162, d166);
	and (d225, d138, d154);
	and (d226, d153, d166);
	and (d227, d144, d150);
	not (d228, d24);
	xor (d229, d170, d177);
	not (d230, d94);
	xor (d231, d118, d145);
	xnor (d232, d158, d161);
	and (d233, d162, d170);
	nor (d234, d160, d173);
	and (d235, d123, d171);
	not (d236, d110);
	not (d237, d16);
	xnor (d238, d153);
	and (d239, d130, d163);
	buf (d240, d143);
	nor (d241, d131, d176);
	buf (d242, d109);
	xnor (d243, d125, d156);
	xnor (d244, d157, d161);
	nor (d245, d122, d125);
	and (d246, d122, d159);
	or (d247, d164, d172);
	or (d248, d139, d162);
	xnor (d249, d171, d176);
	xnor (d250, d157, d169);
	buf (d251, d74);
	xor (d252, d232, d242);
	nor (d253, d202, d205);
	xnor (d254, d184, d202);
	xnor (d255, d201, d210);
	not (d256, d209);
	nor (d257, d237, d242);
	not (d258, d113);
	xor (d259, d207, d214);
	and (d260, d181, d238);
	or (d261, d217, d232);
	xor (d262, d226, d249);
	nand (d263, d194, d220);
	or (d264, d209, d240);
	buf (d265, d12);
	and (d266, d210, d237);
	not (d267, d153);
	buf (d268, d3);
	buf (d269, d100);
	and (d270, d226, d233);
	or (d271, d195, d231);
	xnor (d272, d205, d232);
	xnor (d273, d193, d231);
	nor (d274, d183, d203);
	nor (d275, d205, d218);
	and (d276, d199, d211);
	xor (d277, d188, d215);
	nand (d278, d195, d251);
	or (d279, d202, d223);
	buf (d280, d9);
	or (d281, d223, d226);
	buf (d282, d117);
	and (d283, d195, d217);
	and (d284, d189, d212);
	nor (d285, d203, d231);
	and (d286, d204, d233);
	nand (d287, d188, d215);
	buf (d288, d54);
	nand (d289, d221, d233);
	xnor (d290, d189, d205);
	nand (d291, d213, d214);
	xor (d292, d183, d195);
	and (d293, d190, d199);
	buf (d294, d11);
	xnor (d295, d196, d199);
	nor (d296, d198, d211);
	buf (d297, d249);
	or (d298, d191, d222);
	and (d299, d189, d190);
	xor (d300, d223, d229);
	or (d301, d203, d226);
	buf (d302, d165);
	nand (d303, d181, d206);
	xor (d304, d201, d224);
	xor (d305, d226, d240);
	and (d306, d218, d223);
	buf (d307, d196);
	nor (d308, d181, d190);
	xor (d309, d220, d237);
	buf (d310, d242);
	and (d311, d203, d229);
	buf (d312, d38);
	nor (d313, d201, d230);
	nor (d314, d202, d250);
	buf (d315, d221);
	nor (d316, d184, d240);
	or (d317, d207, d220);
	nor (d318, d192, d213);
	nor (d319, d205, d212);
	not (d320, d134);
	and (d321, d207, d226);
	xor (d322, d230, d239);
	or (d323, d202, d245);
	xnor (d324, d203, d208);
	xor (d325, d199, d249);
	and (d326, d190, d239);
	nand (d327, d201, d228);
	and (d328, d254, d277);
	xor (d329, d269, d292);
	and (d330, d255, d294);
	nand (d331, d286, d312);
	nand (d332, d270, d272);
	nand (d333, d296, d301);
	buf (d334, d323);
	nor (d335, d253, d311);
	xnor (d336, d305, d307);
	nand (d337, d271, d313);
	nor (d338, d255, d327);
	not (d339, d179);
	or (d340, d310, d324);
	nor (d341, d253, d296);
	buf (d342, d276);
	xor (d343, d255, d327);
	not (d344, d138);
	not (d345, d177);
	xor (d346, d335, d338);
	xnor (d347, d332, d335);
	or (d348, d330, d332);
	and (d349, d329, d333);
	nand (d350, d330, d337);
	nor (d351, d329, d336);
	nand (d352, d329, d330);
	nor (d353, d341, d345);
	not (d354, d92);
	and (d355, d341, d344);
	and (d356, d331, d344);
	assign f1 = d354;
	assign f2 = d348;
	assign f3 = d356;
	assign f4 = d355;
endmodule
