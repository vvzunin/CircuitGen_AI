module CCGRCG72( x0, x1, x2, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17, f18, f19 );

	input x0, x1, x2;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17, f18, f19;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314, d315, d316, d317, d318, d319, d320, d321, d322, d323, d324, d325, d326, d327, d328, d329, d330, d331, d332, d333, d334, d335, d336, d337, d338, d339, d340, d341, d342, d343, d344, d345, d346, d347, d348, d349, d350, d351, d352, d353, d354, d355, d356, d357, d358, d359, d360, d361, d362, d363, d364, d365, d366, d367, d368;

	not (d1, x2);
	nor (d2, x0);
	nand (d3, x1, x2);
	nand (d4, x0, x1);
	or (d5, x1, x2);
	nand (d6, x1, x2);
	and (d7, x1, x2);
	nand (d8, x1);
	and (d9, x0, x2);
	nor (d10, x0, x2);
	and (d11, x1, x2);
	buf (d12, x0);
	xor (d13, x1, x2);
	buf (d14, x1);
	nand (d15, x0, x2);
	or (d16, x0, x2);
	nor (d17, x0, x1);
	xnor (d18, x1);
	and (d19, x2);
	not (d20, d13);
	xor (d21, d7, d14);
	xnor (d22, d1, d2);
	not (d23, d19);
	and (d24, d10, d14);
	and (d25, d8, d12);
	nor (d26, d3, d9);
	and (d27, d2, d6);
	xor (d28, d3, d9);
	xnor (d29, d4, d8);
	xor (d30, d6, d15);
	or (d31, d12, d13);
	xor (d32, d15, d19);
	or (d33, d1, d19);
	xor (d34, d7, d12);
	buf (d35, d4);
	nor (d36, d3, d14);
	xnor (d37, d5, d10);
	xor (d38, d8, d14);
	nor (d39, d8, d17);
	or (d40, d11, d12);
	nand (d41, d3, d10);
	nand (d42, d9, d17);
	and (d43, d7, d10);
	not (d44, d8);
	xnor (d45, d10, d18);
	and (d46, d9, d12);
	nand (d47, d7, d19);
	buf (d48, d7);
	and (d49, d10, d14);
	and (d50, d2, d3);
	and (d51, d11, d14);
	xnor (d52, d5, d19);
	nand (d53, d8, d18);
	nand (d54, d5, d15);
	and (d55, d12, d19);
	nand (d56, d13, d19);
	nor (d57, d7, d17);
	nand (d58, d3, d9);
	nor (d59, d1, d13);
	nor (d60, d15, d16);
	xnor (d61, d5, d7);
	not (d62, d42);
	xnor (d63, d27, d55);
	nor (d64, d30, d38);
	xnor (d65, d27, d57);
	buf (d66, d45);
	xor (d67, d31, d51);
	not (d68, d11);
	or (d69, d24, d49);
	xnor (d70, d50, d60);
	nand (d71, d36, d54);
	nor (d72, d30, d52);
	buf (d73, d46);
	or (d74, d36, d44);
	or (d75, d27, d28);
	nand (d76, d27, d42);
	buf (d77, d23);
	nor (d78, d45, d53);
	xnor (d79, d40, d56);
	buf (d80, d24);
	xnor (d81, d35, d49);
	nor (d82, d43, d47);
	xor (d83, d56, d59);
	nor (d84, d48, d61);
	xor (d85, d33, d41);
	and (d86, d22, d52);
	and (d87, d29, d41);
	or (d88, d28, d59);
	xor (d89, d20, d28);
	not (d90, d39);
	and (d91, d43, d61);
	or (d92, d47, d50);
	nor (d93, d46, d52);
	xnor (d94, d58);
	nand (d95, d22, d57);
	not (d96, d27);
	or (d97, d27, d58);
	not (d98, d15);
	and (d99, d34, d36);
	xnor (d100, d49, d56);
	nand (d101, d44, d60);
	nor (d102, d22, d26);
	and (d103, d45, d52);
	not (d104, d32);
	nand (d105, d36, d39);
	xnor (d106, d34, d56);
	or (d107, d36, d37);
	nand (d108, d30, d33);
	buf (d109, d12);
	not (d110, d5);
	xnor (d111, d52, d55);
	xnor (d112, d46, d57);
	nor (d113, d28, d38);
	or (d114, d77, d111);
	or (d115, d72, d106);
	nor (d116, d83, d95);
	not (d117, d23);
	xor (d118, d69, d85);
	xor (d119, d98, d109);
	or (d120, d69, d97);
	xor (d121, d97, d106);
	buf (d122, d80);
	buf (d123, d49);
	nand (d124, d67, d84);
	buf (d125, d73);
	nand (d126, d106, d111);
	xnor (d127, d86, d100);
	nand (d128, d67, d83);
	not (d129, d83);
	nor (d130, d67, d83);
	not (d131, d48);
	buf (d132, d107);
	xor (d133, d71, d74);
	xor (d134, d108);
	buf (d135, d35);
	xor (d136, d74, d93);
	xnor (d137, d71, d91);
	xnor (d138, d85, d111);
	nand (d139, d87, d106);
	not (d140, d44);
	xnor (d141, d117, d132);
	not (d142, d47);
	xor (d143, d119, d121);
	not (d144, d68);
	or (d145, d116, d137);
	xor (d146, d120, d122);
	xor (d147, d133, d138);
	nor (d148, d118, d126);
	xnor (d149, d118, d128);
	not (d150, d10);
	buf (d151, d57);
	and (d152, d129, d138);
	and (d153, d133, d136);
	xor (d154, d117, d130);
	xor (d155, d130, d139);
	buf (d156, d133);
	xnor (d157, d124, d131);
	xnor (d158, d118, d121);
	nor (d159, d127, d135);
	or (d160, d131, d139);
	or (d161, d125, d126);
	xnor (d162, d119, d128);
	nor (d163, d118, d127);
	xor (d164, d118, d128);
	xor (d165, d121, d138);
	nand (d166, d119, d138);
	not (d167, d109);
	not (d168, d24);
	not (d169, d88);
	xnor (d170, d115, d121);
	buf (d171, d112);
	not (d172, d135);
	xnor (d173, d119, d138);
	or (d174, d116, d125);
	buf (d175, d37);
	or (d176, d116, d118);
	xnor (d177, d119, d135);
	not (d178, d45);
	nor (d179, d120, d123);
	nor (d180, d123, d136);
	buf (d181, d40);
	or (d182, d126, d137);
	not (d183, d87);
	and (d184, d118, d133);
	xnor (d185, d117, d130);
	and (d186, d123, d131);
	and (d187, d119, d124);
	not (d188, d56);
	xnor (d189, d133, d138);
	not (d190, d138);
	buf (d191, d116);
	xor (d192, d127, d136);
	nand (d193, d129, d133);
	not (d194, d49);
	nand (d195, d130, d136);
	nor (d196, d119, d122);
	buf (d197, d127);
	or (d198, d118, d122);
	not (d199, d126);
	not (d200, d93);
	and (d201, d116, d130);
	or (d202, d121, d134);
	xnor (d203, d114, d123);
	not (d204, d73);
	not (d205, d120);
	nand (d206, d122, d126);
	buf (d207, d99);
	buf (d208, x2);
	xnor (d209, d119, d125);
	and (d210, d128, d133);
	and (d211, d137, d139);
	and (d212, d114, d130);
	or (d213, d127, d135);
	nand (d214, d118, d120);
	buf (d215, d6);
	not (d216, d134);
	xor (d217, d196, d211);
	nor (d218, d212, d213);
	or (d219, d154, d201);
	nor (d220, d148, d193);
	xor (d221, d141, d207);
	nand (d222, d195, d210);
	nor (d223, d190, d196);
	xnor (d224, d150, d208);
	buf (d225, d164);
	nor (d226, d141, d194);
	and (d227, d155, d208);
	buf (d228, d5);
	or (d229, d171, d182);
	and (d230, d151, d195);
	xor (d231, d178, d204);
	nor (d232, d154, d179);
	buf (d233, d90);
	and (d234, d189, d197);
	and (d235, d160, d173);
	not (d236, d97);
	or (d237, d151, d201);
	or (d238, d204, d212);
	xor (d239, d141, d166);
	or (d240, d186, d206);
	xor (d241, d154, d162);
	nor (d242, d140, d158);
	and (d243, d146, d168);
	nor (d244, d177, d208);
	nor (d245, d167, d205);
	not (d246, d57);
	or (d247, d157, d212);
	or (d248, d147, d160);
	and (d249, d145, d149);
	not (d250, d159);
	xor (d251, d160, d166);
	or (d252, d206, d212);
	nor (d253, d185, d209);
	buf (d254, d50);
	not (d255, d51);
	nor (d256, d156, d165);
	xnor (d257, d192, d203);
	nor (d258, d149, d154);
	xnor (d259, d144, d154);
	xnor (d260, d169, d184);
	nand (d261, d155, d168);
	xor (d262, d170, d185);
	or (d263, d183, d192);
	nand (d264, d175, d178);
	nand (d265, d168, d194);
	buf (d266, d184);
	xnor (d267, d173, d202);
	buf (d268, d67);
	xor (d269, d154, d186);
	nand (d270, d163, d206);
	nor (d271, d157, d164);
	and (d272, d140, d214);
	xor (d273, d152, d190);
	or (d274, d190, d197);
	not (d275, d187);
	and (d276, d186, d211);
	not (d277, d20);
	nand (d278, d154, d182);
	nand (d279, d166, d210);
	nor (d280, d163, d209);
	nor (d281, d170, d172);
	or (d282, d146, d165);
	not (d283, d81);
	or (d284, d208, d210);
	nand (d285, d182, d196);
	nor (d286, d169, d209);
	and (d287, d158, d163);
	nand (d288, d169, d181);
	nand (d289, d155, d163);
	nor (d290, d169, d203);
	or (d291, d179, d214);
	and (d292, d156, d168);
	xnor (d293, d156, d181);
	and (d294, d171, d179);
	and (d295, d173, d180);
	xor (d296, d165, d204);
	not (d297, d150);
	xnor (d298, d148, d152);
	xor (d299, d145, d210);
	xnor (d300, d160, d199);
	buf (d301, d114);
	buf (d302, d95);
	xor (d303, d165);
	xor (d304, d148, d211);
	or (d305, d277, d299);
	nor (d306, d247, d272);
	xnor (d307, d221, d253);
	nor (d308, d290, d304);
	xnor (d309, d220, d257);
	nor (d310, d218, d240);
	or (d311, d260, d299);
	or (d312, d249, d290);
	not (d313, d290);
	nand (d314, d295, d298);
	or (d315, d276, d298);
	nor (d316, d234, d277);
	nand (d317, d233, d281);
	not (d318, d185);
	or (d319, d277, d292);
	nand (d320, d221, d253);
	buf (d321, d115);
	xnor (d322, d236, d240);
	and (d323, d245, d257);
	nor (d324, d222, d302);
	and (d325, d222, d301);
	xnor (d326, d221, d300);
	buf (d327, d68);
	and (d328, d223, d233);
	xor (d329, d276, d300);
	not (d330, d180);
	or (d331, d240, d280);
	xor (d332, d237, d279);
	buf (d333, d189);
	xor (d334, d227, d230);
	xor (d335, d257, d276);
	xnor (d336, d257, d301);
	buf (d337, d130);
	xor (d338, d291, d302);
	and (d339, d302, d303);
	xnor (d340, d230, d273);
	and (d341, d267, d297);
	or (d342, d286, d297);
	buf (d343, d101);
	nand (d344, d232, d290);
	xnor (d345, d228, d250);
	or (d346, d226, d245);
	or (d347, d232, d242);
	nor (d348, d268, d274);
	and (d349, d274);
	not (d350, d221);
	nand (d351, d261, d282);
	nand (d352, d266, d283);
	buf (d353, d211);
	xnor (d354, d226, d278);
	xnor (d355, d248, d284);
	not (d356, d128);
	and (d357, d235, d272);
	and (d358, d243, d262);
	xor (d359, d268, d291);
	and (d360, d248, d300);
	nor (d361, d294, d296);
	nor (d362, d235, d249);
	and (d363, d239, d240);
	and (d364, d230, d303);
	buf (d365, d84);
	xnor (d366, d318, d337);
	not (d367, d356);
	xnor (d368, d358, d362);
	assign f1 = d368;
	assign f2 = d367;
	assign f3 = d367;
	assign f4 = d367;
	assign f5 = d365;
	assign f6 = d368;
	assign f7 = d365;
	assign f8 = d367;
	assign f9 = d367;
	assign f10 = d368;
	assign f11 = d366;
	assign f12 = d367;
	assign f13 = d368;
	assign f14 = d365;
	assign f15 = d367;
	assign f16 = d365;
	assign f17 = d367;
	assign f18 = d368;
	assign f19 = d365;
endmodule
