module CCGRCG10( x0, x1, f1, f2, f3, f4, f5, f6, f7 );

	input x0, x1;
	output f1, f2, f3, f4, f5, f6, f7;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141;

	xnor (d1, x0, x1);
	nor (d2, x0, x1);
	and (d3, x0, x1);
	nor (d4, x0);
	nor (d5, x0, x1);
	xor (d6, x0, x1);
	nand (d7, x0, x1);
	not (d8, x0);
	and (d9, x0);
	or (d10, x0, x1);
	not (d11, x1);
	xnor (d12, x0, x1);
	xor (d13, x1);
	nor (d14, x1);
	or (d15, x0, x1);
	buf (d16, x0);
	xnor (d17, x0);
	or (d18, d7, d13);
	xnor (d19, d6, d14);
	xnor (d20, d7, d13);
	nor (d21, d1, d2);
	xnor (d22, d8, d9);
	and (d23, d1);
	or (d24, d12, d13);
	xor (d25, d7, d11);
	nand (d26, d14, d17);
	xor (d27, d9, d14);
	buf (d28, d9);
	buf (d29, d10);
	xnor (d30, d6, d11);
	nor (d31, d4, d6);
	buf (d32, d3);
	nor (d33, d8, d12);
	xor (d34, d6, d17);
	xor (d35, d8, d9);
	not (d36, d7);
	nor (d37, d3, d5);
	xnor (d38, d4, d15);
	and (d39, d2, d4);
	not (d40, d9);
	not (d41, d1);
	buf (d42, d4);
	nand (d43, d3, d12);
	nor (d44, d5, d17);
	and (d45, d5, d7);
	nand (d46, d9);
	nor (d47, d3, d10);
	or (d48, d7, d10);
	xor (d49, d11, d17);
	not (d50, d13);
	and (d51, d1, d16);
	and (d52, d8, d15);
	xor (d53, d2, d14);
	or (d54, d1, d7);
	and (d55, d3, d15);
	nand (d56, d8, d14);
	buf (d57, d6);
	or (d58, d15, d17);
	xor (d59, d12);
	xor (d60, d10, d12);
	xor (d61, d5, d16);
	not (d62, d2);
	and (d63, d10, d12);
	and (d64, d5, d15);
	not (d65, d14);
	xnor (d66, d1, d3);
	buf (d67, d5);
	buf (d68, d14);
	or (d69, d2, d15);
	nor (d70, d1, d2);
	xor (d71, d4, d5);
	nand (d72, d2, d15);
	or (d73, d9, d15);
	and (d74, d8, d9);
	nand (d75, d3, d15);
	nor (d76, d2, d8);
	buf (d77, d12);
	nor (d78, d3, d13);
	xor (d79, d16, d17);
	nand (d80, d6, d10);
	xor (d81, d12, d14);
	xor (d82, d6, d10);
	buf (d83, d13);
	xor (d84, d4, d9);
	and (d85, d4, d17);
	and (d86, d9, d12);
	or (d87, d14, d16);
	and (d88, d7, d10);
	xor (d89, d1, d12);
	not (d90, d8);
	xor (d91, d6, d13);
	not (d92, d12);
	or (d93, d13, d15);
	nor (d94, d28);
	nand (d95, d37, d51);
	buf (d96, d89);
	nand (d97, d18, d38);
	and (d98, d65, d87);
	xnor (d99, d63, d82);
	buf (d100, d64);
	xnor (d101, d45, d58);
	xnor (d102, d69, d84);
	and (d103, d27, d36);
	xnor (d104, d40, d76);
	and (d105, d44, d91);
	xnor (d106, d26, d44);
	nand (d107, d56, d62);
	xor (d108, d69, d73);
	and (d109, d41, d83);
	nand (d110, d67, d83);
	buf (d111, d79);
	nand (d112, d31, d67);
	buf (d113, d53);
	xor (d114, d25, d38);
	xor (d115, d28, d48);
	not (d116, d87);
	or (d117, d82, d86);
	nor (d118, d60, d75);
	nor (d119, d62, d74);
	xnor (d120, d61, d69);
	xor (d121, d32, d82);
	and (d122, d57, d63);
	not (d123, d38);
	buf (d124, d11);
	nor (d125, d29, d56);
	not (d126, d76);
	nor (d127, d66, d80);
	buf (d128, d78);
	nor (d129, d26, d80);
	nor (d130, d41, d64);
	nand (d131, d47, d62);
	not (d132, d20);
	xnor (d133, d39, d51);
	xnor (d134, d51, d63);
	nand (d135, d33, d68);
	xor (d136, d43, d91);
	or (d137, d42, d71);
	or (d138, d46, d86);
	and (d139, d25, d92);
	not (d140, d68);
	nand (d141, d50, d82);
	assign f1 = d135;
	assign f2 = d141;
	assign f3 = d131;
	assign f4 = d133;
	assign f5 = d118;
	assign f6 = d136;
	assign f7 = d128;
endmodule
