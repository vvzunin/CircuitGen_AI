module CCGRCG436( x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17, f18, f19, f20, f21, f22, f23, f24, f25, f26 );

	input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17, f18, f19, f20, f21, f22, f23, f24, f25, f26;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314, d315, d316, d317, d318, d319, d320, d321, d322, d323, d324, d325, d326, d327, d328, d329, d330, d331, d332, d333, d334, d335, d336, d337, d338, d339, d340, d341, d342, d343, d344, d345, d346, d347, d348, d349, d350, d351, d352, d353, d354, d355, d356, d357, d358, d359, d360, d361, d362, d363, d364, d365, d366, d367, d368, d369, d370, d371, d372, d373, d374, d375, d376, d377, d378, d379, d380, d381, d382, d383, d384, d385, d386, d387, d388, d389, d390, d391, d392, d393, d394, d395, d396, d397, d398, d399, d400, d401, d402, d403, d404, d405, d406, d407, d408, d409, d410, d411, d412, d413, d414, d415, d416, d417, d418, d419, d420, d421, d422, d423, d424, d425, d426, d427, d428, d429, d430, d431, d432, d433, d434, d435, d436, d437, d438, d439, d440, d441, d442, d443, d444, d445, d446, d447, d448, d449, d450, d451, d452, d453, d454, d455, d456, d457, d458, d459, d460, d461, d462, d463, d464, d465, d466, d467, d468, d469, d470, d471, d472, d473, d474, d475, d476, d477, d478, d479, d480, d481, d482, d483, d484, d485, d486, d487, d488, d489, d490, d491, d492, d493, d494, d495, d496, d497, d498, d499, d500, d501, d502, d503, d504, d505, d506, d507, d508, d509, d510, d511, d512, d513, d514, d515, d516, d517, d518, d519, d520, d521, d522, d523, d524, d525, d526, d527, d528, d529, d530, d531, d532, d533, d534, d535, d536, d537, d538, d539, d540, d541, d542, d543, d544, d545, d546, d547, d548, d549, d550, d551, d552, d553, d554, d555, d556, d557, d558, d559, d560, d561, d562, d563, d564, d565, d566, d567, d568, d569, d570, d571, d572, d573, d574, d575, d576, d577, d578, d579, d580, d581, d582, d583, d584, d585, d586, d587, d588, d589, d590, d591, d592, d593, d594, d595, d596, d597, d598, d599, d600, d601, d602, d603, d604, d605, d606, d607, d608, d609, d610, d611, d612, d613, d614, d615, d616, d617, d618, d619, d620, d621, d622, d623, d624, d625, d626, d627, d628, d629, d630, d631, d632, d633, d634, d635, d636, d637, d638, d639, d640, d641, d642, d643, d644, d645, d646, d647, d648, d649, d650, d651, d652, d653, d654, d655, d656, d657, d658, d659, d660, d661, d662, d663, d664, d665, d666, d667, d668, d669, d670, d671, d672, d673, d674, d675, d676, d677, d678, d679, d680, d681, d682, d683, d684, d685, d686, d687, d688, d689, d690, d691, d692, d693, d694, d695, d696, d697, d698, d699, d700, d701, d702, d703, d704, d705, d706, d707, d708, d709, d710, d711, d712, d713, d714, d715, d716, d717, d718, d719, d720, d721, d722, d723, d724, d725, d726, d727, d728, d729, d730, d731, d732, d733, d734, d735, d736, d737, d738, d739, d740, d741, d742, d743, d744, d745, d746, d747, d748, d749, d750, d751, d752, d753, d754, d755, d756, d757, d758, d759;

	nand ( d1, x1, x14);
	not ( d2, x0);
	and ( d3, x11, x27);
	and ( d4, x1, x18);
	buf ( d5, x4);
	nor ( d6, x17, x28);
	xnor ( d7, x15, x26);
	xor ( d8, x8, x27);
	nor ( d9, x19, x22);
	or ( d10, x16, x28);
	or ( d11, x14, x18);
	and ( d12, x8, x29);
	nor ( d13, x18, x19);
	xnor ( d14, x7, x17);
	nor ( d15, x19, x21);
	not ( d16, x11);
	nand ( d17, x17, x28);
	buf ( d18, x29);
	xnor ( d19, x1, x4);
	not ( d20, x7);
	nand ( d21, x15, x24);
	buf ( d22, x24);
	xnor ( d23, x8, x22);
	xor ( d24, x16, x26);
	or ( d25, x18, x26);
	nor ( d26, x17, x21);
	not ( d27, x28);
	or ( d28, x8, x24);
	xnor ( d29, x3, x14);
	not ( d30, x15);
	or ( d31, x13, x27);
	xor ( d32, x28, x29);
	nor ( d33, x8, x17);
	xor ( d34, x5, x26);
	not ( d35, x20);
	and ( d36, x22, x29);
	buf ( d37, x16);
	nor ( d38, x5, x12);
	not ( d39, x29);
	nor ( d40, x0, x27);
	or ( d41, x6, x23);
	nand ( d42, x18, x25);
	or ( d43, x9, x20);
	nor ( d44, x22, x26);
	or ( d45, x24, x26);
	xor ( d46, x21, x22);
	xnor ( d47, x11, x13);
	nand ( d48, x0, x18);
	or ( d49, x6, x10);
	or ( d50, x0, x11);
	and ( d51, x13, x24);
	and ( d52, x13, x29);
	and ( d53, x19, x20);
	nand ( d54, x11, x28);
	xor ( d55, x0, x4);
	not ( d56, x16);
	or ( d57, x4, x23);
	and ( d58, x2, x12);
	nand ( d59, x10, x29);
	xor ( d60, x12, x15);
	nor ( d61, x1, x4);
	nand ( d62, x19, x29);
	or ( d63, x14, x15);
	buf ( d64, x21);
	and ( d65, x2, x16);
	nor ( d66, x9, x14);
	xor ( d67, d7, d55);
	xor ( d68, d6, d26);
	buf ( d69, x15);
	nand ( d70, d42, d63);
	xor ( d71, d30, d50);
	xor ( d72, d2, d64);
	and ( d73, d11, d31);
	xnor ( d74, d35, d36);
	xor ( d75, d22, d47);
	xor ( d76, d58, d64);
	xnor ( d77, d4, d6);
	buf ( d78, x18);
	nor ( d79, d46, d62);
	not ( d80, x18);
	xnor ( d81, d3, d24);
	buf ( d82, d41);
	nand ( d83, d27, d35);
	xor ( d84, d4, d20);
	or ( d85, d21);
	xnor ( d86, d52, d58);
	or ( d87, d23, d36);
	xor ( d88, d24, d39);
	xor ( d89, d4, d45);
	xor ( d90, d3, d48);
	nor ( d91, d11, d49);
	not ( d92, d19);
	xor ( d93, d20, d58);
	or ( d94, d16, d46);
	nand ( d95, d15, d43);
	nand ( d96, d24, d63);
	not ( d97, x14);
	and ( d98, d5, d15);
	and ( d99, d17, d28);
	buf ( d100, d1);
	xnor ( d101, d19, d40);
	not ( d102, x4);
	xnor ( d103, d15, d65);
	nand ( d104, d17, d55);
	and ( d105, d56, d58);
	nand ( d106, d21, d49);
	not ( d107, d5);
	xor ( d108, d4, d10);
	nand ( d109, d54, d59);
	not ( d110, d29);
	and ( d111, d1, d57);
	xor ( d112, d1, d62);
	nand ( d113, d37, d39);
	xor ( d114, d60, d64);
	or ( d115, d22, d25);
	buf ( d116, d11);
	buf ( d117, d7);
	xor ( d118, d52, d62);
	buf ( d119, d50);
	or ( d120, d32, d64);
	or ( d121, d25, d46);
	nand ( d122, d16, d38);
	xor ( d123, d1, d40);
	xnor ( d124, d27, d50);
	nand ( d125, d56, d59);
	nand ( d126, d4, d56);
	and ( d127, d113, d117);
	and ( d128, d71, d103);
	nand ( d129, d79, d98);
	nor ( d130, d92, d102);
	and ( d131, d98, d103);
	or ( d132, d81, d100);
	not ( d133, d24);
	nor ( d134, d82, d120);
	nand ( d135, d105, d113);
	xnor ( d136, d79, d108);
	buf ( d137, d77);
	not ( d138, d36);
	nand ( d139, d98, d115);
	xor ( d140, d73, d109);
	xnor ( d141, d67, d80);
	buf ( d142, d125);
	nor ( d143, d75, d123);
	xor ( d144, d69, d118);
	nand ( d145, d101, d112);
	nor ( d146, d119, d126);
	or ( d147, d97, d104);
	and ( d148, d97, d110);
	nor ( d149, d72, d78);
	xor ( d150, d79, d113);
	buf ( d151, x7);
	nor ( d152, d96, d118);
	and ( d153, d69, d86);
	xor ( d154, d89, d99);
	and ( d155, d85, d90);
	and ( d156, d67, d75);
	or ( d157, d70, d83);
	not ( d158, d80);
	xor ( d159, d68, d83);
	nor ( d160, d77, d79);
	nand ( d161, d67, d73);
	xnor ( d162, d87, d122);
	not ( d163, d111);
	xnor ( d164, d76, d85);
	nand ( d165, d88, d111);
	xor ( d166, d82, d109);
	xor ( d167, d83, d113);
	nor ( d168, d72, d98);
	xnor ( d169, d73, d110);
	or ( d170, d72, d122);
	xor ( d171, d88, d99);
	xor ( d172, d70, d112);
	or ( d173, d115, d123);
	or ( d174, d81, d113);
	nand ( d175, d93, d101);
	xnor ( d176, d79, d81);
	nor ( d177, d72, d108);
	and ( d178, d83, d118);
	xnor ( d179, d112, d116);
	not ( d180, d54);
	xnor ( d181, d74, d120);
	xnor ( d182, d74, d100);
	xnor ( d183, d67, d114);
	nor ( d184, d93, d106);
	nand ( d185, d94, d96);
	or ( d186, d88, d105);
	and ( d187, d71);
	not ( d188, d18);
	and ( d189, d168, d187);
	not ( d190, d177);
	nand ( d191, d142, d173);
	or ( d192, d176, d180);
	xor ( d193, d147, d182);
	not ( d194, d88);
	nor ( d195, d182, d183);
	not ( d196, d155);
	not ( d197, d31);
	or ( d198, d176, d185);
	nand ( d199, d130, d164);
	xnor ( d200, d140, d178);
	xor ( d201, d178, d184);
	xor ( d202, d139, d165);
	and ( d203, d148, d168);
	buf ( d204, d136);
	xnor ( d205, d132, d180);
	not ( d206, x19);
	nand ( d207, d152, d169);
	nor ( d208, d155, d165);
	xnor ( d209, d137, d172);
	nand ( d210, d157, d178);
	xnor ( d211, d173, d177);
	buf ( d212, x14);
	xnor ( d213, d167, d173);
	or ( d214, d163, d170);
	nand ( d215, d145);
	nand ( d216, d166, d176);
	nand ( d217, d190, d204);
	and ( d218, d190, d207);
	xnor ( d219, d200, d210);
	buf ( d220, d16);
	xor ( d221, d189, d212);
	xnor ( d222, d198, d206);
	or ( d223, d193, d197);
	nand ( d224, d189, d197);
	xor ( d225, d199, d208);
	buf ( d226, d85);
	nand ( d227, d199, d200);
	or ( d228, d193, d196);
	or ( d229, d198, d203);
	xor ( d230, d199, d213);
	and ( d231, d197, d206);
	xor ( d232, d189, d203);
	and ( d233, d188, d197);
	nand ( d234, d191, d192);
	and ( d235, d190, d209);
	and ( d236, d201, d210);
	not ( d237, x3);
	and ( d238, d188, d206);
	xor ( d239, d194, d213);
	xnor ( d240, d194, d199);
	xor ( d241, d204, d209);
	nand ( d242, d196, d206);
	and ( d243, d189, d209);
	nor ( d244, d203, d210);
	xnor ( d245, d193, d198);
	and ( d246, d193, d206);
	buf ( d247, d4);
	or ( d248, d202, d210);
	nor ( d249, d194, d204);
	and ( d250, d188, d201);
	xnor ( d251, d211, d215);
	or ( d252, d191, d192);
	and ( d253, d203, d204);
	nand ( d254, d200, d203);
	buf ( d255, d186);
	not ( d256, d41);
	xnor ( d257, d198, d201);
	not ( d258, d168);
	buf ( d259, d173);
	or ( d260, d199, d206);
	or ( d261, d197, d216);
	xnor ( d262, d192, d207);
	xnor ( d263, d206, d216);
	buf ( d264, d212);
	and ( d265, d198, d202);
	nor ( d266, d197, d205);
	buf ( d267, d31);
	and ( d268, d189, d201);
	buf ( d269, d177);
	buf ( d270, d190);
	and ( d271, d191, d210);
	or ( d272, d199, d213);
	buf ( d273, d152);
	buf ( d274, d196);
	xor ( d275, d189, d201);
	xnor ( d276, d191, d215);
	nor ( d277, d194, d216);
	nand ( d278, d206, d213);
	nor ( d279, d196, d198);
	xor ( d280, d202, d215);
	not ( d281, d52);
	and ( d282, d202);
	nand ( d283, d233, d265);
	and ( d284, d234, d259);
	nor ( d285, d217, d270);
	buf ( d286, d222);
	or ( d287, d225, d240);
	not ( d288, x9);
	xor ( d289, d262, d268);
	xor ( d290, d255, d268);
	and ( d291, d230, d270);
	xnor ( d292, d234, d236);
	nor ( d293, d229, d265);
	buf ( d294, d215);
	nor ( d295, d220, d232);
	nor ( d296, d226, d271);
	or ( d297, d230, d239);
	nor ( d298, d226, d266);
	or ( d299, d262, d274);
	nand ( d300, d227, d247);
	buf ( d301, d274);
	xor ( d302, d225, d257);
	buf ( d303, d59);
	not ( d304, x27);
	or ( d305, d246, d263);
	nor ( d306, d220, d244);
	nand ( d307, d249, d258);
	nand ( d308, d218, d277);
	nand ( d309, d241, d244);
	xnor ( d310, d236, d269);
	nor ( d311, d219, d226);
	nand ( d312, d246, d261);
	or ( d313, d237, d275);
	nor ( d314, d267, d280);
	or ( d315, d231, d257);
	nand ( d316, d236, d240);
	nand ( d317, d274, d276);
	nand ( d318, d251, d278);
	xnor ( d319, d243, d281);
	not ( d320, d237);
	nand ( d321, d224, d261);
	not ( d322, d212);
	xor ( d323, d272, d275);
	nand ( d324, d230, d262);
	xor ( d325, d274, d276);
	not ( d326, d265);
	xnor ( d327, d222, d254);
	nand ( d328, d236, d260);
	nand ( d329, d218, d281);
	xor ( d330, d268, d274);
	nor ( d331, d218, d236);
	xor ( d332, d272, d278);
	and ( d333, d238, d248);
	or ( d334, d269, d276);
	nand ( d335, d232, d272);
	xnor ( d336, d271, d276);
	xor ( d337, d244, d267);
	buf ( d338, d118);
	xor ( d339, d262, d281);
	nand ( d340, d241);
	buf ( d341, d280);
	xor ( d342, d267, d278);
	buf ( d343, d70);
	and ( d344, d246, d259);
	nor ( d345, d237, d270);
	buf ( d346, d143);
	or ( d347, d230, d252);
	xnor ( d348, d290, d331);
	xnor ( d349, d298, d303);
	not ( d350, d170);
	not ( d351, d92);
	xnor ( d352, d284, d339);
	xor ( d353, d285, d317);
	xor ( d354, d284, d333);
	xor ( d355, d322, d339);
	xor ( d356, d297, d322);
	nor ( d357, d302, d325);
	xor ( d358, d325, d332);
	buf ( d359, d149);
	not ( d360, d14);
	xnor ( d361, d286);
	and ( d362, d340, d347);
	xor ( d363, d302, d341);
	and ( d364, d286, d294);
	buf ( d365, d287);
	nand ( d366, d283, d338);
	nand ( d367, d292, d329);
	and ( d368, d303, d317);
	or ( d369, d300, d323);
	and ( d370, d295, d344);
	xor ( d371, d313, d327);
	xor ( d372, d294, d305);
	xor ( d373, d284, d335);
	buf ( d374, d132);
	xor ( d375, d330, d333);
	and ( d376, d285, d314);
	nor ( d377, d290, d321);
	xnor ( d378, d306, d343);
	xnor ( d379, d325, d328);
	nor ( d380, d301, d320);
	or ( d381, d305, d316);
	xor ( d382, d315, d344);
	and ( d383, d283, d324);
	not ( d384, d298);
	not ( d385, d32);
	nand ( d386, d319, d320);
	xnor ( d387, d298);
	xnor ( d388, d318, d329);
	buf ( d389, d175);
	xnor ( d390, d298, d328);
	buf ( d391, d165);
	not ( d392, d76);
	nor ( d393, d305, d324);
	nand ( d394, d291, d302);
	or ( d395, d390);
	nand ( d396, d349, d354);
	nand ( d397, d349, d356);
	or ( d398, d368, d385);
	xor ( d399, d391, d394);
	nand ( d400, d362, d369);
	or ( d401, d349, d357);
	xnor ( d402, d371, d391);
	xnor ( d403, d357, d365);
	or ( d404, d349, d388);
	buf ( d405, d240);
	not ( d406, d15);
	xor ( d407, d351, d374);
	xor ( d408, d390);
	and ( d409, d357, d366);
	xnor ( d410, d353, d372);
	nor ( d411, d358, d368);
	nor ( d412, d377, d393);
	xor ( d413, d379, d388);
	xor ( d414, d349, d352);
	xor ( d415, d366, d376);
	and ( d416, d357, d366);
	nor ( d417, d359, d369);
	not ( d418, d300);
	and ( d419, d376, d382);
	buf ( d420, d22);
	xnor ( d421, d367, d379);
	not ( d422, d69);
	not ( d423, d259);
	and ( d424, d358, d384);
	xor ( d425, d350, d384);
	nor ( d426, d348, d376);
	buf ( d427, d355);
	and ( d428, d361, d364);
	or ( d429, d386, d393);
	nor ( d430, d348, d389);
	and ( d431, d355, d358);
	or ( d432, d392, d394);
	xor ( d433, d350, d392);
	or ( d434, d379);
	or ( d435, d375, d382);
	nor ( d436, d362, d366);
	nor ( d437, d380, d387);
	nand ( d438, d366, d379);
	xor ( d439, d372, d385);
	not ( d440, d356);
	nor ( d441, d378, d392);
	or ( d442, d349, d362);
	nor ( d443, d369, d376);
	and ( d444, d364, d365);
	and ( d445, d363, d380);
	or ( d446, d362, d372);
	or ( d447, d371, d391);
	buf ( d448, d94);
	xor ( d449, d396, d440);
	xor ( d450, d411, d425);
	nand ( d451, d415, d441);
	xnor ( d452, d429, d446);
	nand ( d453, d438, d443);
	not ( d454, d328);
	xor ( d455, d398, d403);
	nand ( d456, d406, d442);
	not ( d457, d204);
	buf ( d458, d144);
	buf ( d459, d271);
	and ( d460, d397, d413);
	xor ( d461, d416, d431);
	nor ( d462, d405, d410);
	and ( d463, d416, d423);
	and ( d464, d440);
	xnor ( d465, d412, d420);
	xnor ( d466, d409, d422);
	and ( d467, d406, d418);
	or ( d468, d401, d424);
	xnor ( d469, d405, d426);
	nand ( d470, d435, d445);
	or ( d471, d422, d428);
	or ( d472, d422, d445);
	nor ( d473, d403, d428);
	not ( d474, d53);
	or ( d475, d395, d402);
	and ( d476, d397, d399);
	nand ( d477, d400, d439);
	not ( d478, d173);
	buf ( d479, d238);
	or ( d480, d401, d441);
	and ( d481, d406, d432);
	or ( d482, d405, d417);
	not ( d483, d355);
	buf ( d484, d39);
	nand ( d485, d395, d420);
	buf ( d486, d375);
	not ( d487, d91);
	xor ( d488, d418, d431);
	xnor ( d489, d406, d442);
	and ( d490, d438, d445);
	xnor ( d491, d404, d420);
	buf ( d492, d192);
	nand ( d493, d406, d445);
	nor ( d494, d430, d437);
	and ( d495, d397, d409);
	xnor ( d496, d422, d430);
	xnor ( d497, d436, d441);
	nor ( d498, d398, d420);
	nand ( d499, d395, d397);
	and ( d500, d411, d437);
	and ( d501, d405, d414);
	nand ( d502, d408, d446);
	not ( d503, d340);
	not ( d504, d427);
	or ( d505, d399, d411);
	nand ( d506, d397);
	nor ( d507, d419, d440);
	nand ( d508, d420, d429);
	xnor ( d509, d397, d419);
	xnor ( d510, d412, d418);
	xor ( d511, d427, d442);
	xnor ( d512, d403, d407);
	or ( d513, d403, d419);
	or ( d514, d437, d438);
	and ( d515, d420, d447);
	xor ( d516, d400, d434);
	not ( d517, d44);
	buf ( d518, d148);
	xnor ( d519, d453, d494);
	buf ( d520, d9);
	and ( d521, d470, d471);
	buf ( d522, d336);
	or ( d523, d486, d489);
	and ( d524, d449, d450);
	nor ( d525, d501, d517);
	xor ( d526, d501, d502);
	xnor ( d527, d457, d458);
	nand ( d528, d468, d490);
	and ( d529, d458, d481);
	and ( d530, d455, d515);
	xnor ( d531, d464, d479);
	nand ( d532, d457, d460);
	nor ( d533, d472, d510);
	nand ( d534, d451, d497);
	nand ( d535, d462, d514);
	and ( d536, d480, d482);
	nor ( d537, d498, d515);
	not ( d538, d207);
	xnor ( d539, d458, d477);
	buf ( d540, d109);
	nor ( d541, d455, d513);
	or ( d542, d461, d493);
	nand ( d543, d448, d516);
	xnor ( d544, d473, d517);
	nand ( d545, d458, d476);
	xnor ( d546, d491, d496);
	or ( d547, d501, d515);
	buf ( d548, d245);
	not ( d549, d374);
	xnor ( d550, d463, d476);
	nor ( d551, d449, d496);
	nand ( d552, d486, d496);
	xnor ( d553, d465, d507);
	buf ( d554, d324);
	or ( d555, d491, d506);
	or ( d556, d477, d497);
	xnor ( d557, d458, d492);
	xnor ( d558, d471, d509);
	xnor ( d559, d484, d492);
	not ( d560, d87);
	xnor ( d561, d495, d507);
	or ( d562, d464, d509);
	or ( d563, d478, d510);
	nor ( d564, d465, d490);
	and ( d565, d498, d514);
	and ( d566, d454, d506);
	xor ( d567, d522, d550);
	or ( d568, d565, d566);
	or ( d569, d568);
	xnor ( d570, d567);
	not ( d571, d511);
	buf ( d572, d241);
	xnor ( d573, d568);
	nor ( d574, d568);
	nor ( d575, d567);
	xor ( d576, d567);
	nor ( d577, d572, d576);
	or ( d578, d572, d574);
	xor ( d579, d574, d576);
	xnor ( d580, d570, d574);
	xor ( d581, d570, d571);
	xor ( d582, d571, d576);
	xnor ( d583, d569, d576);
	xnor ( d584, d573, d574);
	or ( d585, d570, d572);
	buf ( d586, d343);
	nor ( d587, d570, d573);
	xor ( d588, d571, d574);
	and ( d589, d569, d571);
	not ( d590, d351);
	not ( d591, d136);
	buf ( d592, d123);
	xor ( d593, d571, d575);
	and ( d594, d569, d576);
	buf ( d595, d14);
	or ( d596, d569, d576);
	nand ( d597, d569, d574);
	not ( d598, d218);
	buf ( d599, d576);
	nor ( d600, d569, d576);
	and ( d601, d570, d571);
	buf ( d602, d209);
	and ( d603, d574, d575);
	nor ( d604, d572, d573);
	xor ( d605, d573, d575);
	nand ( d606, d572);
	nor ( d607, d575, d576);
	xnor ( d608, d570, d574);
	nor ( d609, d570, d574);
	nor ( d610, d572, d574);
	nor ( d611, d571, d574);
	nand ( d612, d569, d573);
	xor ( d613, d573, d575);
	or ( d614, d574, d576);
	buf ( d615, d277);
	or ( d616, d571, d572);
	xnor ( d617, d573, d575);
	nor ( d618, d571, d576);
	xnor ( d619, d569, d574);
	xnor ( d620, d569, d571);
	xor ( d621, d571, d575);
	not ( d622, d563);
	nand ( d623, d578, d603);
	and ( d624, d577, d610);
	buf ( d625, d316);
	nand ( d626, d594, d619);
	or ( d627, d586, d587);
	buf ( d628, d583);
	nand ( d629, d595, d618);
	and ( d630, d609, d612);
	buf ( d631, d457);
	xor ( d632, d587, d602);
	and ( d633, d596, d607);
	xor ( d634, d601, d620);
	nor ( d635, d593, d614);
	xor ( d636, d586, d608);
	and ( d637, d593, d605);
	nor ( d638, d596, d601);
	and ( d639, d581, d584);
	or ( d640, d583, d590);
	nor ( d641, d594, d610);
	nand ( d642, d601, d608);
	nand ( d643, d578, d580);
	or ( d644, d583, d588);
	not ( d645, d287);
	nor ( d646, d592, d613);
	xor ( d647, d593, d620);
	xnor ( d648, d581, d621);
	buf ( d649, d305);
	not ( d650, d620);
	xor ( d651, d579, d594);
	and ( d652, d600, d619);
	nand ( d653, d578, d598);
	nor ( d654, d583, d610);
	and ( d655, d586, d621);
	nand ( d656, d584, d618);
	or ( d657, d588, d604);
	or ( d658, d582, d588);
	and ( d659, d580, d603);
	nand ( d660, d578, d610);
	xor ( d661, d593, d600);
	not ( d662, d604);
	or ( d663, d579, d617);
	xor ( d664, d586, d601);
	not ( d665, d336);
	nand ( d666, d607, d613);
	buf ( d667, d543);
	or ( d668, d596, d612);
	or ( d669, d588, d618);
	and ( d670, d586, d603);
	buf ( d671, d19);
	not ( d672, d554);
	xnor ( d673, d586, d611);
	and ( d674, d578, d617);
	nor ( d675, d596, d598);
	nor ( d676, d593, d603);
	nor ( d677, d590, d617);
	nand ( d678, d577, d582);
	and ( d679, d595, d602);
	nor ( d680, d582, d609);
	buf ( d681, d337);
	and ( d682, d603, d610);
	buf ( d683, d327);
	and ( d684, d599);
	or ( d685, d591, d614);
	or ( d686, d581, d612);
	and ( d687, d663, d684);
	xnor ( d688, d622, d671);
	or ( d689, d647, d680);
	nand ( d690, d662, d671);
	not ( d691, d302);
	and ( d692, d632, d646);
	nor ( d693, d638, d655);
	nor ( d694, d654);
	nor ( d695, d641, d677);
	nor ( d696, d631, d669);
	and ( d697, d647, d652);
	not ( d698, d668);
	buf ( d699, d294);
	nand ( d700, d660, d661);
	and ( d701, d649, d676);
	or ( d702, d656, d669);
	or ( d703, d646, d650);
	buf ( d704, x10);
	not ( d705, d516);
	and ( d706, d656, d685);
	xnor ( d707, d674, d684);
	or ( d708, d624, d672);
	buf ( d709, d589);
	not ( d710, d249);
	nor ( d711, d623, d637);
	xnor ( d712, d634, d661);
	nor ( d713, d642, d653);
	nor ( d714, d643, d679);
	nor ( d715, d649, d655);
	nor ( d716, d664, d679);
	nand ( d717, d652, d664);
	not ( d718, d500);
	or ( d719, d637, d664);
	nand ( d720, d643, d685);
	buf ( d721, d137);
	or ( d722, d632, d633);
	or ( d723, d659, d670);
	xor ( d724, d653, d670);
	buf ( d725, d369);
	xor ( d726, d646);
	and ( d727, d651, d679);
	or ( d728, d661, d686);
	and ( d729, d646, d672);
	or ( d730, d668, d679);
	xor ( d731, d689, d692);
	xnor ( d732, d697, d713);
	nor ( d733, d716, d729);
	xnor ( d734, d716, d725);
	nor ( d735, d706, d712);
	nand ( d736, d708, d730);
	and ( d737, d701, d717);
	xor ( d738, d706, d729);
	nor ( d739, d687, d715);
	nor ( d740, d687, d714);
	and ( d741, d689, d706);
	not ( d742, d322);
	buf ( d743, x13);
	not ( d744, d722);
	xnor ( d745, d708, d712);
	nand ( d746, d696, d707);
	xnor ( d747, d699, d702);
	nor ( d748, d700, d714);
	nand ( d749, d706, d715);
	xnor ( d750, d717, d719);
	xnor ( d751, d700, d714);
	or ( d752, d691, d724);
	and ( d753, d688, d722);
	nor ( d754, d689, d700);
	xor ( d755, d690, d696);
	xnor ( d756, d710, d722);
	xor ( d757, d691, d713);
	buf ( d758, d742);
	buf ( d759, d76);
	assign f1 = d759;
	assign f2 = d759;
	assign f3 = d759;
	assign f4 = d759;
	assign f5 = d759;
	assign f6 = d759;
	assign f7 = d759;
	assign f8 = d758;
	assign f9 = d758;
	assign f10 = d758;
	assign f11 = d758;
	assign f12 = d759;
	assign f13 = d758;
	assign f14 = d759;
	assign f15 = d759;
	assign f16 = d758;
	assign f17 = d758;
	assign f18 = d758;
	assign f19 = d758;
	assign f20 = d758;
	assign f21 = d759;
	assign f22 = d759;
	assign f23 = d758;
	assign f24 = d759;
	assign f25 = d758;
	assign f26 = d758;
endmodule
