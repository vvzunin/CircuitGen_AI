module CCGRCG4( x0, x1, f1, f2, f3, f4 );

	input x0, x1;
	output f1, f2, f3, f4;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314, d315, d316, d317, d318, d319, d320, d321, d322, d323, d324, d325, d326, d327, d328, d329, d330, d331, d332, d333, d334, d335, d336, d337, d338, d339, d340, d341, d342, d343, d344, d345, d346, d347, d348, d349, d350, d351, d352, d353, d354, d355, d356, d357, d358, d359, d360, d361, d362, d363, d364, d365, d366, d367, d368, d369, d370, d371, d372, d373, d374, d375, d376, d377, d378, d379, d380, d381, d382, d383, d384, d385, d386, d387, d388, d389, d390, d391, d392, d393, d394, d395, d396, d397, d398, d399, d400, d401, d402, d403, d404, d405, d406, d407, d408, d409, d410, d411, d412, d413, d414, d415, d416, d417, d418, d419, d420, d421, d422, d423, d424, d425, d426, d427, d428, d429, d430, d431, d432, d433;

	xor (d1, x0, x1);
	xor (d2, x0, x1);
	nor (d3, x0);
	nand (d4, x0);
	buf (d5, x0);
	and (d6, x0, x1);
	nand (d7, x1);
	or (d8, x0);
	not (d9, x0);
	nand (d10, x0, x1);
	nor (d11, x1);
	xnor (d12, x0, x1);
	nor (d13, x0, x1);
	buf (d14, x1);
	nand (d15, d3, d13);
	xnor (d16, d5);
	xor (d17, d4, d12);
	and (d18, d9, d11);
	or (d19, d3, d6);
	nand (d20, d2, d11);
	and (d21, d8, d11);
	or (d22, d10);
	not (d23, d2);
	xnor (d24, d7, d13);
	and (d25, d5, d11);
	xor (d26, d1, d8);
	xor (d27, d5, d14);
	nand (d28, d2, d5);
	nor (d29, d3, d7);
	and (d30, d2, d5);
	nand (d31, d8, d9);
	nor (d32, d2, d4);
	or (d33, d11, d14);
	xor (d34, d5, d7);
	or (d35, d5, d13);
	or (d36, d6, d8);
	or (d37, d7, d10);
	nand (d38, d11, d13);
	buf (d39, d12);
	and (d40, d3, d13);
	not (d41, d4);
	buf (d42, d3);
	xnor (d43, d10, d11);
	nand (d44, d10, d11);
	not (d45, d9);
	xnor (d46, d3, d6);
	buf (d47, d5);
	and (d48, d5, d14);
	and (d49, d4, d11);
	xor (d50, d4, d7);
	xnor (d51, d8, d13);
	nor (d52, d1, d10);
	and (d53, d11, d13);
	xor (d54, d1, d4);
	xnor (d55, d3, d7);
	nor (d56, d1, d4);
	buf (d57, d4);
	xor (d58, d14);
	nor (d59, d1, d3);
	nor (d60, d2, d5);
	nor (d61, d47, d57);
	not (d62, d39);
	buf (d63, d22);
	xnor (d64, d28, d57);
	nor (d65, d31, d46);
	and (d66, d23, d40);
	buf (d67, d36);
	nor (d68, d50, d54);
	nand (d69, d39, d43);
	and (d70, d29, d41);
	nand (d71, d36, d37);
	or (d72, d16, d19);
	and (d73, d28, d51);
	nand (d74, d17, d45);
	and (d75, d27, d33);
	and (d76, d16, d19);
	xor (d77, d19);
	xor (d78, d23, d43);
	not (d79, d27);
	xor (d80, d15, d18);
	nor (d81, d27, d46);
	or (d82, d24, d40);
	not (d83, d29);
	xnor (d84, d37, d54);
	buf (d85, d21);
	not (d86, d41);
	nor (d87, d43, d47);
	nor (d88, d26, d39);
	nand (d89, d39, d48);
	and (d90, d21, d29);
	xor (d91, d35, d44);
	or (d92, d33, d59);
	and (d93, d27, d30);
	not (d94, d54);
	nand (d95, d20, d24);
	nand (d96, d45, d55);
	not (d97, d48);
	xor (d98, d45, d46);
	not (d99, d17);
	or (d100, d31, d38);
	and (d101, d24, d38);
	nor (d102, d17, d24);
	xor (d103, d28, d42);
	and (d104, d31, d58);
	buf (d105, d26);
	nor (d106, d18, d37);
	not (d107, d10);
	xnor (d108, d54);
	or (d109, d22, d59);
	xnor (d110, d16, d47);
	xor (d111, d20, d54);
	and (d112, d29, d47);
	not (d113, d57);
	or (d114, d30, d39);
	xor (d115, d26, d56);
	xnor (d116, d20, d44);
	not (d117, d42);
	nor (d118, d18, d42);
	not (d119, d47);
	or (d120, d24, d41);
	nand (d121, d39, d41);
	not (d122, d43);
	nand (d123, d34, d41);
	or (d124, d18, d19);
	or (d125, d32, d53);
	buf (d126, d52);
	xnor (d127, d43);
	and (d128, d15, d20);
	or (d129, d15, d27);
	not (d130, d13);
	and (d131, d18, d29);
	or (d132, d24, d47);
	not (d133, d18);
	xnor (d134, d24, d26);
	xnor (d135, d16, d37);
	nor (d136, d30, d48);
	xnor (d137, d27, d55);
	xor (d138, d46, d50);
	buf (d139, d45);
	buf (d140, d57);
	xor (d141, d27, d58);
	xnor (d142, d49, d57);
	nor (d143, d48, d49);
	and (d144, d31, d46);
	not (d145, d56);
	xor (d146, d21, d31);
	and (d147, d50, d57);
	nor (d148, d47, d48);
	nand (d149, d15, d16);
	nor (d150, d32, d46);
	not (d151, d12);
	xor (d152, d48, d51);
	and (d153, d66, d144);
	or (d154, d83, d149);
	and (d155, d113, d128);
	or (d156, d70, d142);
	nor (d157, d66, d98);
	nand (d158, d83, d132);
	xnor (d159, d73, d150);
	xnor (d160, d74, d139);
	and (d161, d155, d159);
	nand (d162, d153, d157);
	nand (d163, d154, d160);
	not (d164, d138);
	nor (d165, d157, d159);
	nand (d166, d153, d158);
	or (d167, d156, d160);
	xnor (d168, d158, d160);
	nand (d169, d153, d155);
	and (d170, d157, d159);
	nand (d171, d153, d156);
	nand (d172, d154, d158);
	or (d173, d153, d156);
	nor (d174, d156, d159);
	or (d175, d153, d157);
	xor (d176, d153, d156);
	nor (d177, d153, d154);
	nand (d178, d153, d155);
	nor (d179, d153, d155);
	nor (d180, d155, d158);
	xor (d181, d157, d160);
	not (d182, d140);
	not (d183, d128);
	buf (d184, d63);
	not (d185, d103);
	xor (d186, d158, d160);
	and (d187, d153, d156);
	or (d188, d154, d160);
	xnor (d189, d157, d158);
	or (d190, d154, d158);
	xor (d191, d156, d157);
	xnor (d192, d159, d160);
	and (d193, d154, d156);
	xnor (d194, d153, d158);
	xor (d195, d157, d158);
	or (d196, d159);
	xor (d197, d155, d159);
	or (d198, d156, d159);
	xnor (d199, d158, d160);
	and (d200, d153, d159);
	xor (d201, d153, d155);
	xor (d202, d155, d156);
	buf (d203, d40);
	not (d204, d153);
	and (d205, d155, d157);
	xnor (d206, d154, d160);
	xnor (d207, d153, d157);
	nand (d208, d154, d157);
	and (d209, d153, d159);
	nor (d210, d155, d158);
	and (d211, d158, d160);
	buf (d212, d117);
	not (d213, d99);
	or (d214, d155);
	nand (d215, d157, d159);
	or (d216, d156);
	nand (d217, d153, d160);
	or (d218, d156, d160);
	nor (d219, d156);
	xor (d220, d159, d160);
	and (d221, d169, d170);
	xnor (d222, d185);
	buf (d223, d13);
	not (d224, d184);
	not (d225, d159);
	or (d226, d177, d207);
	nand (d227, d165, d167);
	xor (d228, d212, d214);
	nand (d229, d178, d181);
	and (d230, d168, d171);
	buf (d231, d11);
	or (d232, d193, d212);
	xor (d233, d163, d185);
	not (d234, d181);
	and (d235, d179, d188);
	xnor (d236, d187, d203);
	xor (d237, d193, d215);
	and (d238, d175, d186);
	or (d239, d175, d179);
	or (d240, d176, d178);
	and (d241, d162, d173);
	xnor (d242, d194, d197);
	nand (d243, d168, d203);
	xnor (d244, d191, d192);
	or (d245, d162, d173);
	and (d246, d177, d184);
	or (d247, d188, d218);
	nor (d248, d174, d200);
	not (d249, d143);
	buf (d250, d167);
	or (d251, d175, d190);
	or (d252, d164, d174);
	nand (d253, d174, d210);
	nand (d254, d172, d198);
	xnor (d255, d172, d203);
	buf (d256, d50);
	and (d257, d212, d217);
	buf (d258, d89);
	xor (d259, d187, d209);
	buf (d260, d215);
	nor (d261, d204, d220);
	not (d262, d11);
	xnor (d263, d176, d198);
	and (d264, d175, d215);
	xor (d265, d177, d220);
	or (d266, d166, d180);
	nand (d267, d190, d219);
	not (d268, d178);
	xor (d269, d163, d203);
	xnor (d270, d245, d268);
	xnor (d271, d241, d242);
	buf (d272, d104);
	buf (d273, d239);
	not (d274, d154);
	or (d275, d256, d263);
	buf (d276, d252);
	not (d277, d90);
	nor (d278, d234, d262);
	and (d279, d224, d267);
	xor (d280, d221, d260);
	or (d281, d229, d268);
	nor (d282, d229, d240);
	nand (d283, d225);
	nor (d284, d228, d240);
	buf (d285, d139);
	xnor (d286, d239, d243);
	nand (d287, d229, d238);
	not (d288, d219);
	and (d289, d255, d258);
	xor (d290, d236, d261);
	or (d291, d244, d255);
	and (d292, d221, d263);
	nor (d293, d246, d260);
	nand (d294, d247, d260);
	xnor (d295, d241, d258);
	nand (d296, d235, d258);
	nor (d297, d226, d241);
	not (d298, d226);
	xor (d299, d240, d267);
	not (d300, d185);
	nor (d301, d244, d263);
	nand (d302, d222, d247);
	xor (d303, d229, d242);
	nor (d304, d224, d236);
	nor (d305, d241, d243);
	and (d306, d251, d266);
	nand (d307, d224, d232);
	xor (d308, d223, d241);
	nand (d309, d226, d237);
	buf (d310, d90);
	and (d311, d243, d260);
	not (d312, d105);
	not (d313, d75);
	xnor (d314, d222, d259);
	nand (d315, d225, d256);
	not (d316, d264);
	nand (d317, d233, d238);
	xnor (d318, d261, d268);
	and (d319, d233, d243);
	nor (d320, d225, d269);
	nor (d321, d253, d257);
	and (d322, d222, d250);
	not (d323, d91);
	buf (d324, d241);
	xnor (d325, d227, d233);
	nand (d326, d256, d263);
	xor (d327, d223, d226);
	xnor (d328, d223, d269);
	or (d329, d237, d249);
	xnor (d330, d227, d263);
	nor (d331, d224, d261);
	or (d332, d222, d231);
	or (d333, d238, d252);
	xor (d334, d253, d264);
	and (d335, d222, d267);
	and (d336, d223, d266);
	buf (d337, d246);
	xor (d338, d251, d262);
	xnor (d339, d226, d235);
	and (d340, d317, d319);
	buf (d341, d222);
	xnor (d342, d282, d324);
	or (d343, d300, d315);
	not (d344, d192);
	not (d345, d203);
	and (d346, d274, d330);
	xnor (d347, d303, d321);
	buf (d348, d161);
	xnor (d349, d309, d313);
	or (d350, d294, d312);
	xor (d351, d281, d326);
	or (d352, d274, d281);
	nand (d353, d291, d329);
	nor (d354, d278, d294);
	nor (d355, d289, d311);
	or (d356, d298, d303);
	or (d357, d292, d316);
	xnor (d358, d302, d327);
	xor (d359, d307, d325);
	nand (d360, d275, d319);
	or (d361, d275, d312);
	nand (d362, d289, d293);
	or (d363, d299, d316);
	xnor (d364, d277, d324);
	nand (d365, d298);
	xor (d366, d275, d336);
	xor (d367, d286, d325);
	xor (d368, d270, d298);
	buf (d369, d43);
	xnor (d370, d278, d315);
	or (d371, d284, d294);
	nor (d372, d312, d333);
	xnor (d373, d327, d331);
	not (d374, d195);
	buf (d375, d262);
	or (d376, d274, d304);
	buf (d377, d68);
	xnor (d378, d306, d331);
	and (d379, d297, d299);
	buf (d380, d71);
	and (d381, d296, d312);
	nor (d382, d277, d326);
	and (d383, d274, d328);
	xor (d384, d325, d329);
	nor (d385, d275, d318);
	buf (d386, d334);
	nor (d387, d284, d319);
	not (d388, d122);
	nand (d389, d294, d333);
	xor (d390, d311, d335);
	xnor (d391, d281, d292);
	not (d392, d217);
	xor (d393, d273, d308);
	and (d394, d279, d300);
	xor (d395, d280, d307);
	buf (d396, d268);
	buf (d397, d230);
	and (d398, d307, d335);
	nor (d399, d306, d324);
	xor (d400, d307, d315);
	xnor (d401, d275, d304);
	not (d402, d130);
	nand (d403, d309, d313);
	xnor (d404, d302, d335);
	xor (d405, d291, d302);
	nand (d406, d355, d383);
	or (d407, d364, d381);
	or (d408, d341, d371);
	buf (d409, d176);
	or (d410, d349, d384);
	and (d411, d350, d358);
	xor (d412, d371, d374);
	buf (d413, d295);
	nor (d414, d344, d378);
	buf (d415, d405);
	and (d416, d347, d396);
	and (d417, d362, d378);
	nand (d418, d381, d387);
	and (d419, d351, d403);
	not (d420, d293);
	nor (d421, d363, d380);
	or (d422, d379, d381);
	buf (d423, d309);
	xnor (d424, d369, d391);
	and (d425, d341, d347);
	nor (d426, d347, d365);
	and (d427, d346, d363);
	nor (d428, d368, d370);
	or (d429, d343, d357);
	buf (d430, d190);
	xor (d431, d394, d399);
	nand (d432, d377, d384);
	nand (d433, d379, d393);
	assign f1 = d426;
	assign f2 = d420;
	assign f3 = d428;
	assign f4 = d425;
endmodule
