module CCGRCG106( x0, x1, x2, x3, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17 );

	input x0, x1, x2, x3;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314, d315, d316, d317, d318, d319, d320, d321, d322, d323, d324, d325, d326, d327, d328, d329, d330, d331, d332, d333, d334, d335, d336, d337, d338, d339, d340, d341, d342, d343, d344, d345, d346, d347, d348, d349, d350, d351, d352, d353, d354, d355, d356, d357, d358, d359, d360, d361, d362, d363, d364, d365, d366, d367, d368, d369, d370, d371, d372, d373, d374, d375, d376, d377, d378, d379, d380, d381, d382, d383, d384, d385, d386, d387, d388, d389;

	xor (d1, x0, x1);
	buf (d2, x0);
	nor (d3, x0, x3);
	buf (d4, x3);
	or (d5, x0, x1);
	or (d6, x0, x1);
	xor (d7, x1);
	or (d8, x1, x2);
	nand (d9, x0, x1);
	xor (d10, x0, x1);
	xnor (d11, x1, x3);
	nor (d12, x0, x3);
	xnor (d13, x0, x3);
	or (d14, x3);
	xor (d15, x1, x3);
	nand (d16, x2, x3);
	xor (d17, x0, x3);
	nand (d18, x1, x3);
	xnor (d19, x1, x2);
	xnor (d20, x2);
	nor (d21, x3);
	nor (d22, x0, x1);
	or (d23, x0, x2);
	nor (d24, x1, x3);
	nor (d25, x0, x2);
	nand (d26, x0, x2);
	nand (d27, x1, x2);
	or (d28, x0, x2);
	and (d29, x1, x3);
	nand (d30, x1, x3);
	not (d31, x2);
	not (d32, x0);
	xnor (d33, x2, x3);
	xnor (d34, x3);
	nor (d35, x1, x2);
	nor (d36, x2);
	and (d37, x0, x2);
	xnor (d38, x0, x1);
	xnor (d39, x1, x3);
	and (d40, x0, x1);
	and (d41, x1, x3);
	nand (d42, x2);
	or (d43, x0, x3);
	nor (d44, x2, x3);
	buf (d45, x1);
	or (d46, x2);
	not (d47, x1);
	xor (d48, x1, x2);
	and (d49, x1, x2);
	xnor (d50, x1);
	or (d51, x1, x2);
	xnor (d52, x0, x1);
	xor (d53, x2, x3);
	nor (d54, x1);
	nand (d55, x0, x3);
	nand (d56, x1, x2);
	nor (d57, x1, x2);
	nand (d58, x0, x3);
	xnor (d59, x0);
	or (d60, x0, x3);
	nor (d61, x0, x1);
	nor (d62, x0);
	xor (d63, x2);
	and (d64, x0);
	buf (d65, x2);
	and (d66, d1, d58);
	not (d67, d6);
	nor (d68, d60, d61);
	and (d69, d4, d44);
	xor (d70, d5, d50);
	and (d71, d41, d55);
	nor (d72, d24, d29);
	nor (d73, d16, d30);
	not (d74, d60);
	buf (d75, d65);
	not (d76, d62);
	or (d77, d16, d29);
	xor (d78, d18, d33);
	nand (d79, d23, d63);
	nor (d80, d2, d39);
	not (d81, d43);
	buf (d82, d26);
	xnor (d83, d17, d19);
	nor (d84, d26, d31);
	nand (d85, d16, d62);
	not (d86, d3);
	nor (d87, d33, d39);
	xnor (d88, d31, d39);
	buf (d89, d32);
	nand (d90, d1, d16);
	xor (d91, d17, d42);
	xor (d92, d6, d22);
	nor (d93, d3, d25);
	xor (d94, d10, d62);
	or (d95, d55, d57);
	and (d96, d10, d12);
	and (d97, d38, d54);
	not (d98, d9);
	nand (d99, d4, d5);
	xor (d100, d57, d58);
	and (d101, d2, d36);
	xor (d102, d12, d32);
	buf (d103, d8);
	xor (d104, d17, d36);
	and (d105, d23, d61);
	and (d106, d31, d34);
	or (d107, d35, d64);
	buf (d108, d53);
	or (d109, d26, d51);
	nor (d110, d10, d18);
	xor (d111, d36, d55);
	xnor (d112, d9, d58);
	buf (d113, d61);
	or (d114, d35, d45);
	and (d115, d15, d35);
	not (d116, d50);
	buf (d117, d33);
	xor (d118, d7);
	nand (d119, d10, d34);
	or (d120, d7, d25);
	xnor (d121, d1, d25);
	xor (d122, d11, d45);
	xnor (d123, d5, d19);
	xnor (d124, d45, d57);
	xnor (d125, d42, d64);
	or (d126, d59, d63);
	not (d127, d24);
	xnor (d128, d14, d53);
	xnor (d129, d4, d64);
	nor (d130, d17, d34);
	xnor (d131, d29, d34);
	and (d132, d6, d34);
	not (d133, d47);
	and (d134, d50, d64);
	xnor (d135, d9, d31);
	nor (d136, d46, d49);
	xor (d137, d14, d43);
	buf (d138, d40);
	nor (d139, d14, d47);
	or (d140, d3, d18);
	and (d141, d36, d45);
	nor (d142, d53, d55);
	nand (d143, d51, d54);
	not (d144, d40);
	buf (d145, d59);
	nand (d146, d47, d57);
	or (d147, d1, d32);
	or (d148, d29, d45);
	buf (d149, d28);
	or (d150, d25, d52);
	and (d151, d58, d60);
	xor (d152, d48, d60);
	xnor (d153, d58, d59);
	nor (d154, d3, d62);
	buf (d155, d88);
	not (d156, d72);
	or (d157, d95, d120);
	nand (d158, d97);
	and (d159, d81, d151);
	xor (d160, d119, d148);
	xor (d161, d83, d90);
	and (d162, d68, d152);
	nor (d163, d88, d138);
	not (d164, d120);
	nor (d165, d69, d113);
	or (d166, d74, d87);
	nand (d167, d103, d138);
	buf (d168, d55);
	or (d169, d100, d112);
	nand (d170, d77, d96);
	nand (d171, d85, d134);
	not (d172, d39);
	buf (d173, d60);
	xor (d174, d86, d116);
	nand (d175, d94, d118);
	xor (d176, d100, d128);
	or (d177, d90, d127);
	nand (d178, d134, d139);
	xor (d179, d67, d99);
	nor (d180, d105, d112);
	buf (d181, d44);
	or (d182, d134, d137);
	and (d183, d92, d124);
	buf (d184, d15);
	or (d185, d66, d122);
	nor (d186, d78, d135);
	xor (d187, d135, d139);
	xor (d188, d108, d149);
	not (d189, d100);
	xnor (d190, d96, d127);
	nand (d191, d106, d110);
	xnor (d192, d97, d145);
	and (d193, d77, d108);
	xnor (d194, d72, d116);
	xnor (d195, d69, d81);
	or (d196, d141, d154);
	xnor (d197, d104, d131);
	xor (d198, d103, d138);
	xor (d199, d79, d113);
	or (d200, d84, d140);
	buf (d201, d34);
	or (d202, d102, d152);
	xnor (d203, d83, d120);
	nor (d204, d81, d83);
	buf (d205, d107);
	nor (d206, d99, d116);
	or (d207, d72, d147);
	not (d208, d154);
	xor (d209, d75, d131);
	buf (d210, d121);
	xnor (d211, d96, d112);
	and (d212, d108, d114);
	or (d213, d92, d103);
	buf (d214, d75);
	nand (d215, d113, d150);
	buf (d216, d17);
	nor (d217, d127, d137);
	buf (d218, d142);
	nor (d219, d66, d108);
	nor (d220, d98, d104);
	xor (d221, d189, d215);
	xor (d222, d192, d216);
	buf (d223, d4);
	xnor (d224, d182, d191);
	nand (d225, d156, d160);
	xor (d226, d223, d224);
	nor (d227, d223, d224);
	not (d228, d140);
	nand (d229, d222, d223);
	or (d230, d221, d223);
	or (d231, d223, d224);
	and (d232, d222, d224);
	nor (d233, d222);
	xor (d234, d221, d222);
	buf (d235, d116);
	and (d236, d221, d224);
	xor (d237, d223, d225);
	nor (d238, d223);
	or (d239, d224, d225);
	nand (d240, d223, d225);
	nand (d241, d223, d224);
	and (d242, d222, d225);
	xor (d243, d224, d225);
	nor (d244, d221, d223);
	xnor (d245, d223, d224);
	or (d246, d222, d224);
	nand (d247, d223, d225);
	or (d248, d221, d224);
	xnor (d249, d221, d223);
	xnor (d250, d224);
	xor (d251, d224, d225);
	nand (d252, d224, d225);
	xnor (d253, d221, d223);
	xnor (d254, d222, d224);
	xnor (d255, d223, d225);
	or (d256, d223, d224);
	nor (d257, d225);
	nor (d258, d222, d225);
	or (d259, d223, d225);
	buf (d260, d42);
	xnor (d261, d223, d225);
	nor (d262, d222, d224);
	buf (d263, d106);
	xor (d264, d221);
	xnor (d265, d224, d225);
	nor (d266, d221, d225);
	nor (d267, d222, d225);
	xnor (d268, d223, d224);
	not (d269, d1);
	nor (d270, d221, d222);
	and (d271, d221, d224);
	nand (d272, d221, d225);
	and (d273, d222, d223);
	and (d274, d224, d225);
	nor (d275, d223, d225);
	not (d276, d77);
	and (d277, d223, d224);
	nand (d278, d222, d224);
	nor (d279, d221, d224);
	not (d280, d92);
	not (d281, d22);
	nor (d282, d223, d225);
	nor (d283, d224, d225);
	or (d284, d221, d222);
	not (d285, x3);
	xnor (d286, d224, d225);
	xor (d287, d222, d223);
	xnor (d288, d221, d225);
	xor (d289, d223);
	or (d290, d221, d223);
	xnor (d291, d221, d224);
	nand (d292, d223);
	nor (d293, d222, d223);
	buf (d294, d202);
	or (d295, d221);
	buf (d296, d169);
	xor (d297, d221, d223);
	or (d298, d223);
	xnor (d299, d221);
	and (d300, d221, d222);
	or (d301, d222, d223);
	nand (d302, d238, d239);
	and (d303, d244, d295);
	xnor (d304, d236, d291);
	xnor (d305, d262, d287);
	buf (d306, d127);
	nand (d307, d230, d242);
	and (d308, d244, d297);
	nand (d309, d260, d297);
	buf (d310, d251);
	or (d311, d276, d299);
	and (d312, d271, d284);
	nor (d313, d299, d301);
	nand (d314, d239, d278);
	xor (d315, d230, d287);
	buf (d316, d139);
	not (d317, d83);
	buf (d318, d36);
	xor (d319, d268, d288);
	nand (d320, d260, d263);
	xnor (d321, d238, d243);
	xnor (d322, d237, d275);
	nand (d323, d281, d288);
	xnor (d324, d245);
	nor (d325, d233, d281);
	or (d326, d233, d268);
	xor (d327, d259, d273);
	not (d328, d213);
	xnor (d329, d270, d278);
	buf (d330, d73);
	nand (d331, d241, d293);
	not (d332, d68);
	nor (d333, d251, d268);
	or (d334, d240, d250);
	nor (d335, d228, d280);
	or (d336, d264, d266);
	xor (d337, d255, d270);
	buf (d338, d293);
	xor (d339, d230, d281);
	xor (d340, d242, d286);
	not (d341, d8);
	or (d342, d272, d296);
	not (d343, d182);
	xnor (d344, d268, d300);
	or (d345, d265, d301);
	xnor (d346, d231, d284);
	buf (d347, d284);
	xnor (d348, d250, d263);
	buf (d349, d173);
	not (d350, d261);
	buf (d351, d152);
	and (d352, d226, d280);
	nor (d353, d231, d291);
	or (d354, d269, d297);
	not (d355, d162);
	nand (d356, d236, d244);
	not (d357, d143);
	nand (d358, d245, d286);
	not (d359, d202);
	nand (d360, d247, d260);
	and (d361, d261, d295);
	or (d362, d254, d293);
	nand (d363, d267, d300);
	buf (d364, d51);
	nor (d365, d227, d242);
	or (d366, d228, d256);
	xor (d367, d247, d251);
	nor (d368, d230, d237);
	xnor (d369, d294, d296);
	nor (d370, d280, d294);
	and (d371, d236, d277);
	buf (d372, d237);
	not (d373, d220);
	buf (d374, d39);
	nor (d375, d261, d293);
	not (d376, d66);
	buf (d377, d46);
	or (d378, d292, d301);
	and (d379, d230, d247);
	xnor (d380, d233, d300);
	nand (d381, d289, d292);
	nand (d382, d232, d247);
	xnor (d383, d244, d246);
	and (d384, d228, d298);
	xnor (d385, d238, d284);
	buf (d386, d134);
	nor (d387, d282, d289);
	not (d388, d25);
	xnor (d389, d227, d280);
	assign f1 = d352;
	assign f2 = d313;
	assign f3 = d302;
	assign f4 = d372;
	assign f5 = d312;
	assign f6 = d358;
	assign f7 = d320;
	assign f8 = d336;
	assign f9 = d348;
	assign f10 = d347;
	assign f11 = d311;
	assign f12 = d325;
	assign f13 = d318;
	assign f14 = d378;
	assign f15 = d354;
	assign f16 = d374;
	assign f17 = d373;
endmodule
