module CCGRCG18( x0, x1, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11 );

	input x0, x1;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208;

	buf (d1, x0);
	xor (d2, x0);
	not (d3, x1);
	xnor (d4, x0, x1);
	or (d5, x0, x1);
	and (d6, x0);
	or (d7, x0, x1);
	and (d8, x0, x1);
	nor (d9, x0);
	nand (d10, x0, x1);
	xnor (d11, x1);
	xor (d12, x0, x1);
	nor (d13, x0, x1);
	xnor (d14, x0);
	xor (d15, x0, x1);
	nor (d16, x0, x1);
	or (d17, x1);
	buf (d18, x1);
	nand (d19, x1);
	nand (d20, x0, x1);
	xor (d21, x1);
	or (d22, x0);
	not (d23, x0);
	and (d24, x1);
	nor (d25, x1);
	and (d26, x0, x1);
	not (d27, d12);
	and (d28, d10, d23);
	buf (d29, d6);
	xnor (d30, d17, d22);
	and (d31, d10, d17);
	nor (d32, d16, d19);
	xnor (d33, d2, d5);
	xor (d34, d11);
	nor (d35, d17, d22);
	and (d36, d18, d22);
	and (d37, d8, d21);
	and (d38, d22, d23);
	or (d39, d16, d21);
	not (d40, d6);
	nor (d41, d12, d17);
	or (d42, d1, d21);
	nor (d43, d15, d16);
	xor (d44, d6, d17);
	and (d45, d13, d21);
	and (d46, d17, d26);
	xnor (d47, d10, d21);
	not (d48, d17);
	xor (d49, d19, d23);
	nand (d50, d15, d17);
	nand (d51, d4, d24);
	buf (d52, d3);
	xnor (d53, d3, d16);
	nor (d54, d6, d24);
	xor (d55, d8, d23);
	or (d56, d9, d16);
	and (d57, d3, d20);
	nand (d58, d3, d17);
	or (d59, d6, d24);
	and (d60, d14, d18);
	xor (d61, d9, d12);
	nor (d62, d2, d21);
	nor (d63, d21, d25);
	xor (d64, d4, d14);
	and (d65, d1, d4);
	xor (d66, d3, d15);
	not (d67, d18);
	buf (d68, d23);
	not (d69, d15);
	or (d70, d2, d21);
	nor (d71, d8, d20);
	xnor (d72, d16, d22);
	or (d73, d27, d42);
	xor (d74, d48, d58);
	nor (d75, d73);
	not (d76, d54);
	not (d77, d44);
	or (d78, d73, d74);
	not (d79, d69);
	and (d80, d73, d74);
	nor (d81, d73, d74);
	or (d82, d74);
	not (d83, d16);
	nor (d84, d74);
	xor (d85, d73, d74);
	xnor (d86, d74);
	or (d87, d73);
	and (d88, d74);
	xor (d89, d73, d74);
	not (d90, d10);
	buf (d91, d18);
	nor (d92, d73, d74);
	not (d93, d25);
	buf (d94, d64);
	xnor (d95, d73, d74);
	nand (d96, d73, d74);
	not (d97, d62);
	buf (d98, d69);
	nand (d99, d73, d74);
	buf (d100, d38);
	and (d101, d73);
	nand (d102, d73);
	not (d103, d29);
	not (d104, d4);
	and (d105, d73, d74);
	xnor (d106, d73);
	not (d107, d5);
	not (d108, d40);
	xor (d109, d73);
	xor (d110, d74);
	buf (d111, d4);
	nand (d112, d87, d91);
	xnor (d113, d77, d79);
	not (d114, d87);
	nand (d115, d93, d109);
	xor (d116, d100, d111);
	or (d117, d80, d90);
	nand (d118, d82, d91);
	and (d119, d96, d99);
	and (d120, d79, d83);
	or (d121, d76, d83);
	or (d122, d82, d87);
	or (d123, d80, d110);
	nor (d124, d80, d83);
	nor (d125, d114, d115);
	not (d126, d47);
	xnor (d127, d112, d116);
	nor (d128, d119, d124);
	nor (d129, d113, d116);
	and (d130, d117, d120);
	nand (d131, d113, d115);
	nand (d132, d115, d118);
	xor (d133, d120, d124);
	nor (d134, d122);
	or (d135, d116, d123);
	buf (d136, d68);
	or (d137, d112, d115);
	buf (d138, d11);
	not (d139, d92);
	nor (d140, d123, d124);
	buf (d141, d85);
	buf (d142, d73);
	xnor (d143, d119, d122);
	and (d144, d115, d118);
	xor (d145, d117, d118);
	and (d146, d112, d117);
	and (d147, d117, d124);
	not (d148, d94);
	xnor (d149, d134, d140);
	not (d150, d96);
	not (d151, d19);
	and (d152, d143, d148);
	or (d153, d136, d147);
	or (d154, d128, d132);
	and (d155, d144, d145);
	nand (d156, d129, d137);
	xor (d157, d125, d130);
	nand (d158, d139, d143);
	xnor (d159, d139, d146);
	buf (d160, d144);
	nand (d161, d126, d142);
	xnor (d162, d126, d148);
	xor (d163, d126, d139);
	xnor (d164, d137, d139);
	buf (d165, d35);
	or (d166, d125, d143);
	not (d167, d108);
	nor (d168, d141, d145);
	xor (d169, d141, d143);
	nand (d170, d131, d141);
	xnor (d171, d148);
	xor (d172, d133, d143);
	nand (d173, d136, d145);
	not (d174, d53);
	nand (d175, d131, d133);
	xnor (d176, d127, d131);
	nor (d177, d127, d137);
	xnor (d178, d135, d140);
	not (d179, d129);
	or (d180, d129, d132);
	or (d181, d130, d135);
	nand (d182, d132, d145);
	xnor (d183, d130, d136);
	nor (d184, d130, d148);
	not (d185, d132);
	nor (d186, d132, d140);
	or (d187, d136, d146);
	nor (d188, d129, d134);
	xor (d189, d127, d128);
	xor (d190, d129, d141);
	buf (d191, d37);
	buf (d192, d62);
	not (d193, d3);
	xnor (d194, d129, d138);
	not (d195, d28);
	buf (d196, d19);
	xnor (d197, d139, d140);
	xnor (d198, d125, d131);
	nor (d199, d132, d142);
	and (d200, d125, d140);
	nor (d201, d136, d141);
	buf (d202, d41);
	nand (d203, d140, d146);
	and (d204, d142, d148);
	nor (d205, d129, d137);
	xor (d206, d128, d141);
	nor (d207, d131, d133);
	buf (d208, d63);
	assign f1 = d164;
	assign f2 = d173;
	assign f3 = d167;
	assign f4 = d154;
	assign f5 = d167;
	assign f6 = d154;
	assign f7 = d191;
	assign f8 = d168;
	assign f9 = d198;
	assign f10 = d149;
	assign f11 = d163;
endmodule
