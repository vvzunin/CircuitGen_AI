module CCGRCG188( x0, x1, x2, x3, x4, x5, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17, f18, f19, f20 );

	input x0, x1, x2, x3, x4, x5;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17, f18, f19, f20;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294;

	xnor (d1, x3, x4);
	buf (d2, x5);
	xor (d3, x2, x4);
	and (d4, x3);
	buf (d5, x2);
	xor (d6, x0, x4);
	xor (d7, x0, x3);
	or (d8, x3, x5);
	not (d9, x2);
	nand (d10, x0, x2);
	or (d11, x1, x4);
	buf (d12, x3);
	and (d13, x1, x3);
	xor (d14, x1, x2);
	or (d15, x2, x4);
	not (d16, x3);
	not (d17, x4);
	nor (d18, x2, x4);
	not (d19, x5);
	and (d20, x2, x3);
	or (d21, x0, x3);
	xnor (d22, x1);
	nand (d23, x0, x3);
	or (d24, x1);
	xor (d25, x2, x5);
	and (d26, x3, x5);
	nor (d27, x1, x2);
	or (d28, x1, x4);
	xor (d29, x0, x4);
	not (d30, x1);
	or (d31, x5);
	xor (d32, x4, x5);
	xnor (d33, x1, x5);
	xnor (d34, x2, x5);
	buf (d35, x0);
	or (d36, x1, x5);
	xnor (d37, x0, x1);
	xnor (d38, x0, x2);
	nor (d39, x2, x4);
	or (d40, x4, x5);
	nand (d41, x2);
	or (d42, x2, x3);
	nor (d43, x2, x3);
	nor (d44, x3);
	nand (d45, x1, x5);
	not (d46, x0);
	xnor (d47, x0, x4);
	xnor (d48, x0, x5);
	nor (d49, x0, x2);
	and (d50, x0, x2);
	and (d51, x3, x4);
	or (d52, x3, x4);
	buf (d53, x4);
	xor (d54, x3);
	xnor (d55, x2, x4);
	and (d56, x1, x5);
	or (d57, x1, x2);
	nor (d58, x4, x5);
	and (d59, x0, x4);
	nor (d60, x4, x5);
	xnor (d61, x0, x4);
	or (d62, d18, d26);
	nor (d63, d10, d52);
	xor (d64, d45, d46);
	nor (d65, d29, d44);
	or (d66, d7, d59);
	or (d67, d12, d19);
	buf (d68, d3);
	xor (d69, d27, d31);
	buf (d70, d50);
	nand (d71, d5, d45);
	xnor (d72, d4, d49);
	nand (d73, d2, d12);
	not (d74, d25);
	not (d75, d59);
	not (d76, d7);
	buf (d77, d32);
	nand (d78, d4, d48);
	or (d79, d3, d29);
	buf (d80, d42);
	and (d81, d9, d20);
	not (d82, d30);
	nor (d83, d1, d44);
	buf (d84, d23);
	not (d85, d49);
	xnor (d86, d11, d33);
	or (d87, d39, d54);
	nor (d88, d4, d43);
	or (d89, d38, d43);
	buf (d90, d4);
	nand (d91, d12, d28);
	nand (d92, d31, d39);
	buf (d93, d49);
	nor (d94, d36, d54);
	nor (d95, d24, d39);
	xnor (d96, d27, d31);
	or (d97, d8, d12);
	nor (d98, d34, d60);
	buf (d99, d31);
	xor (d100, d40, d44);
	xor (d101, d12, d18);
	nand (d102, d33, d53);
	not (d103, d46);
	or (d104, d9, d12);
	nor (d105, d38, d54);
	or (d106, d11, d58);
	buf (d107, d34);
	and (d108, d13, d57);
	xnor (d109, d11, d22);
	or (d110, d3, d35);
	nor (d111, d33, d47);
	nor (d112, d16, d31);
	xor (d113, d56, d58);
	nor (d114, d1, d45);
	nand (d115, d41, d60);
	and (d116, d22, d26);
	nand (d117, d27, d33);
	xnor (d118, d19, d38);
	nand (d119, d14, d26);
	nand (d120, d30, d53);
	or (d121, d1, d55);
	xnor (d122, d5, d9);
	nand (d123, d23, d35);
	and (d124, d23, d42);
	not (d125, d14);
	and (d126, d16, d53);
	or (d127, d41, d42);
	xnor (d128, d48, d50);
	nor (d129, d8, d48);
	or (d130, d27, d49);
	nand (d131, d6, d24);
	or (d132, d5, d29);
	xor (d133, d3, d33);
	nor (d134, d31, d43);
	xnor (d135, d12, d32);
	xor (d136, d23, d46);
	xnor (d137, d3, d25);
	xor (d138, d41, d53);
	nand (d139, d9, d21);
	nand (d140, d11);
	xor (d141, d1, d15);
	xor (d142, d28, d38);
	or (d143, d15, d36);
	nor (d144, d6, d48);
	xnor (d145, d41, d61);
	not (d146, d15);
	xor (d147, d20, d58);
	buf (d148, d13);
	nor (d149, d11, d14);
	xnor (d150, d3, d50);
	xnor (d151, d18, d32);
	buf (d152, d38);
	and (d153, d16, d59);
	buf (d154, d83);
	buf (d155, d150);
	buf (d156, d82);
	or (d157, d154, d155);
	not (d158, d6);
	xnor (d159, d154, d155);
	nand (d160, d154, d155);
	nor (d161, d159, d160);
	and (d162, d156, d159);
	not (d163, d40);
	nor (d164, d160);
	xor (d165, d157, d160);
	nand (d166, d157, d158);
	or (d167, d156);
	nand (d168, d156);
	and (d169, d157, d158);
	not (d170, d144);
	or (d171, d157);
	nor (d172, d157, d160);
	xnor (d173, d157, d158);
	nor (d174, d159);
	and (d175, d158, d159);
	not (d176, d124);
	not (d177, d95);
	nor (d178, d157, d159);
	or (d179, d157, d160);
	xor (d180, d156, d160);
	not (d181, d29);
	buf (d182, d159);
	or (d183, d158, d159);
	xor (d184, d159);
	xnor (d185, d159, d160);
	xnor (d186, d158, d160);
	buf (d187, d72);
	and (d188, d159);
	xor (d189, d157);
	xor (d190, d156, d160);
	not (d191, d39);
	not (d192, d136);
	xor (d193, d156, d159);
	buf (d194, d104);
	and (d195, d157);
	or (d196, d157, d159);
	nand (d197, d159, d160);
	buf (d198, d94);
	nand (d199, d160);
	nor (d200, d158, d159);
	xor (d201, d156, d157);
	xor (d202, d158, d159);
	and (d203, d171, d175);
	xor (d204, d166, d201);
	xor (d205, d171, d202);
	not (d206, d42);
	nand (d207, d171, d194);
	not (d208, d100);
	xnor (d209, d192, d193);
	nor (d210, d190, d201);
	not (d211, d77);
	not (d212, d99);
	xor (d213, d209, d210);
	or (d214, d204, d207);
	xnor (d215, d207);
	buf (d216, d197);
	nor (d217, d205, d210);
	xor (d218, d207, d210);
	nor (d219, d205, d209);
	nor (d220, d206, d211);
	and (d221, d204, d211);
	or (d222, d210);
	nand (d223, d204, d210);
	buf (d224, d77);
	not (d225, d27);
	buf (d226, d185);
	not (d227, d184);
	or (d228, d207, d211);
	or (d229, d205, d206);
	nor (d230, d205);
	buf (d231, d60);
	nand (d232, d204, d208);
	xnor (d233, d205, d207);
	nand (d234, d204, d209);
	xor (d235, d204, d205);
	xor (d236, d223, d230);
	buf (d237, d43);
	buf (d238, d208);
	and (d239, d225, d234);
	buf (d240, d89);
	nand (d241, d213, d215);
	nand (d242, d212, d218);
	buf (d243, d193);
	nand (d244, d218, d219);
	xnor (d245, d212, d223);
	nand (d246, d222, d223);
	xnor (d247, d218, d227);
	nor (d248, d216, d227);
	nand (d249, d220, d228);
	buf (d250, d199);
	xnor (d251, d212, d215);
	xor (d252, d218, d222);
	nor (d253, d215, d235);
	nor (d254, d218, d233);
	nor (d255, d222, d234);
	nor (d256, d219, d229);
	and (d257, d219, d234);
	xnor (d258, d212, d227);
	not (d259, d37);
	buf (d260, d22);
	not (d261, d61);
	nor (d262, d252, d254);
	not (d263, d16);
	nand (d264, d242, d250);
	xnor (d265, d241, d256);
	not (d266, d80);
	nand (d267, d242, d249);
	xor (d268, d237, d241);
	not (d269, d13);
	xnor (d270, d236, d241);
	xor (d271, d252, d257);
	buf (d272, d184);
	nor (d273, d252, d255);
	and (d274, d243, d254);
	xnor (d275, d247, d257);
	nand (d276, d237, d244);
	and (d277, d239, d254);
	and (d278, d245, d253);
	and (d279, d249, d258);
	xor (d280, d253);
	xor (d281, d241, d244);
	nor (d282, d237, d240);
	xor (d283, d252, d253);
	buf (d284, d221);
	buf (d285, d175);
	or (d286, d268, d281);
	or (d287, d271, d281);
	nand (d288, d275, d281);
	not (d289, d143);
	nor (d290, d270, d276);
	xor (d291, d265, d270);
	not (d292, d91);
	xor (d293, d271, d281);
	not (d294, d85);
	assign f1 = d292;
	assign f2 = d293;
	assign f3 = d290;
	assign f4 = d284;
	assign f5 = d286;
	assign f6 = d290;
	assign f7 = d290;
	assign f8 = d288;
	assign f9 = d286;
	assign f10 = d289;
	assign f11 = d287;
	assign f12 = d291;
	assign f13 = d285;
	assign f14 = d288;
	assign f15 = d290;
	assign f16 = d294;
	assign f17 = d287;
	assign f18 = d290;
	assign f19 = d291;
	assign f20 = d288;
endmodule
