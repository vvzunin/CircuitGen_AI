module CCGRCG2( x0, x1, f1, f2 );

	input x0, x1;
	output f1, f2;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295;

	not (d1, x1);
	or (d2, x1);
	xnor (d3, x1);
	buf (d4, x0);
	nand (d5, x1);
	or (d6, x0, x1);
	nor (d7, x0, x1);
	nand (d8, x0);
	nor (d9, x0, x1);
	and (d10, x1);
	not (d11, x0);
	nand (d12, x0, x1);
	or (d13, x0, x1);
	xnor (d14, x0, x1);
	xnor (d15, d8, d13);
	or (d16, d4, d9);
	xor (d17, d1, d3);
	nand (d18, d6, d13);
	nor (d19, d10, d12);
	or (d20, d2, d8);
	xnor (d21, d6, d9);
	nor (d22, d9, d11);
	nand (d23, d7, d9);
	nand (d24, d4, d11);
	not (d25, d12);
	buf (d26, d13);
	xnor (d27, d2, d10);
	xor (d28, d10, d12);
	xnor (d29, d2, d6);
	not (d30, d4);
	nand (d31, d5, d7);
	xnor (d32, d7);
	buf (d33, d3);
	nand (d34, d3, d4);
	xnor (d35, d8, d9);
	nand (d36, d1, d3);
	or (d37, d10, d14);
	xor (d38, d5, d13);
	buf (d39, d4);
	not (d40, d2);
	nand (d41, d9, d13);
	xor (d42, d2, d14);
	and (d43, d2, d8);
	not (d44, d8);
	nor (d45, d1, d11);
	nor (d46, d1, d2);
	xor (d47, d10, d13);
	and (d48, d6, d8);
	xor (d49, d2, d8);
	nand (d50, d10, d13);
	or (d51, d4, d10);
	xnor (d52, d2, d10);
	and (d53, d5, d14);
	xor (d54, d4, d6);
	xnor (d55, d11, d13);
	or (d56, d8, d9);
	xor (d57, d2, d7);
	buf (d58, d10);
	or (d59, d1, d14);
	and (d60, d3, d9);
	xnor (d61, d2, d14);
	and (d62, d7, d13);
	xnor (d63, d7, d10);
	buf (d64, d6);
	and (d65, d5, d13);
	and (d66, d5, d14);
	xor (d67, d9, d11);
	not (d68, d9);
	and (d69, d7, d10);
	and (d70, d1, d6);
	xor (d71, d3, d4);
	not (d72, d3);
	not (d73, d6);
	buf (d74, d1);
	and (d75, d2, d5);
	or (d76, d4, d8);
	not (d77, d1);
	xor (d78, d2, d13);
	xor (d79, d4, d13);
	and (d80, d2, d7);
	nand (d81, d6, d14);
	and (d82, d1, d11);
	buf (d83, d8);
	buf (d84, d5);
	xnor (d85, d39, d57);
	nand (d86, d26, d40);
	nand (d87, d35, d39);
	or (d88, d64, d76);
	nand (d89, d38, d50);
	nand (d90, d33, d36);
	nor (d91, d48, d52);
	nand (d92, d49, d82);
	not (d93, d75);
	xor (d94, d26, d54);
	or (d95, d69, d79);
	nor (d96, d20, d71);
	buf (d97, d18);
	xnor (d98, d44, d70);
	and (d99, d22, d81);
	buf (d100, d11);
	xnor (d101, d15, d58);
	nand (d102, d16, d48);
	nor (d103, d34, d68);
	nor (d104, d15, d40);
	or (d105, d36, d38);
	nor (d106, d61, d84);
	not (d107, d52);
	xnor (d108, d61, d67);
	xor (d109, d19, d23);
	and (d110, d29, d73);
	buf (d111, d64);
	and (d112, d24, d41);
	and (d113, d30, d44);
	nand (d114, d55, d75);
	not (d115, d54);
	or (d116, d60, d73);
	and (d117, d18, d31);
	xnor (d118, d19, d57);
	nor (d119, d48, d65);
	not (d120, d65);
	nor (d121, d36, d68);
	not (d122, d41);
	not (d123, d66);
	and (d124, d18, d77);
	xnor (d125, d15, d29);
	or (d126, d42, d79);
	not (d127, d74);
	and (d128, d17, d61);
	not (d129, d40);
	nor (d130, d39, d81);
	xor (d131, d36, d42);
	buf (d132, d42);
	xor (d133, d40, d59);
	and (d134, d61, d74);
	or (d135, d25, d71);
	xnor (d136, d35, d81);
	nor (d137, d19, d74);
	buf (d138, d50);
	nor (d139, d34, d78);
	buf (d140, d68);
	buf (d141, d22);
	xnor (d142, d24, d62);
	or (d143, d29, d77);
	or (d144, d53, d60);
	nor (d145, d44, d75);
	buf (d146, d40);
	xor (d147, d16, d57);
	or (d148, d15, d78);
	xnor (d149, d30, d57);
	xor (d150, d38, d83);
	or (d151, d34, d38);
	nor (d152, d56, d70);
	and (d153, d21, d40);
	nand (d154, d24, d54);
	xor (d155, d59, d72);
	nor (d156, d16, d21);
	not (d157, d17);
	not (d158, d64);
	or (d159, d24, d37);
	nand (d160, d40, d45);
	or (d161, d102, d116);
	not (d162, d94);
	not (d163, d136);
	not (d164, d157);
	buf (d165, d28);
	xor (d166, d97, d142);
	or (d167, d102, d155);
	nor (d168, d89, d159);
	buf (d169, d80);
	nor (d170, d134, d145);
	and (d171, d136, d146);
	nand (d172, d90, d103);
	not (d173, d104);
	not (d174, d158);
	and (d175, d135, d136);
	xnor (d176, d102, d122);
	not (d177, d118);
	xnor (d178, d143, d150);
	and (d179, d86, d132);
	xor (d180, d111, d138);
	nand (d181, d109, d156);
	not (d182, d61);
	xnor (d183, d165, d166);
	xor (d184, d174, d179);
	and (d185, d163, d179);
	xor (d186, d172, d173);
	nand (d187, d166, d180);
	xor (d188, d165, d177);
	xor (d189, d161, d163);
	nand (d190, d166, d168);
	nand (d191, d163, d167);
	or (d192, d167, d177);
	buf (d193, d158);
	not (d194, d53);
	nor (d195, d168, d173);
	and (d196, d163, d168);
	and (d197, d179, d180);
	or (d198, d179);
	nor (d199, d169, d175);
	buf (d200, d99);
	not (d201, d128);
	not (d202, d139);
	xor (d203, d165, d173);
	xnor (d204, d165, d178);
	xnor (d205, d162);
	xor (d206, d172, d181);
	and (d207, d170, d180);
	and (d208, d168, d176);
	not (d209, d174);
	nor (d210, d164, d175);
	and (d211, d166, d172);
	buf (d212, x1);
	nand (d213, d169, d170);
	or (d214, d161, d176);
	and (d215, d163, d176);
	or (d216, d174, d180);
	and (d217, d170, d176);
	xnor (d218, d165, d175);
	nand (d219, d171, d177);
	and (d220, d169, d178);
	and (d221, d166, d177);
	buf (d222, d2);
	or (d223, d163, d176);
	or (d224, d172, d177);
	not (d225, d114);
	xor (d226, d165, d170);
	not (d227, d55);
	and (d228, d164, d166);
	not (d229, d121);
	xnor (d230, d175, d181);
	or (d231, d163, d181);
	or (d232, d168, d170);
	xnor (d233, d169, d182);
	xor (d234, d167, d175);
	xor (d235, d168, d180);
	and (d236, d174, d180);
	xnor (d237, d165, d172);
	buf (d238, d100);
	xor (d239, d210);
	or (d240, d224, d226);
	nand (d241, d194, d196);
	and (d242, d190, d231);
	nor (d243, d184, d192);
	buf (d244, d229);
	xnor (d245, d191, d227);
	and (d246, d190, d236);
	xor (d247, d191, d222);
	or (d248, d194, d228);
	nand (d249, d188, d203);
	not (d250, d15);
	or (d251, d203, d238);
	or (d252, d218, d224);
	nor (d253, d183, d202);
	nor (d254, d203, d224);
	xnor (d255, d223, d234);
	not (d256, d219);
	not (d257, d16);
	nor (d258, d210, d215);
	or (d259, d186, d191);
	buf (d260, d143);
	nor (d261, d228, d238);
	or (d262, d200, d212);
	not (d263, d207);
	xnor (d264, d201, d212);
	not (d265, d39);
	or (d266, d185, d202);
	nand (d267, d189, d220);
	buf (d268, d41);
	xnor (d269, d209, d234);
	xor (d270, d224, d230);
	nand (d271, d216, d234);
	xor (d272, d210, d230);
	xor (d273, d218, d230);
	nand (d274, d188, d221);
	xnor (d275, d196, d238);
	xor (d276, d193, d232);
	or (d277, d211, d212);
	xor (d278, d196, d221);
	and (d279, d195, d228);
	buf (d280, d209);
	buf (d281, d144);
	xor (d282, d251, d274);
	or (d283, d261, d264);
	nor (d284, d255, d271);
	xnor (d285, d268, d278);
	or (d286, d258, d270);
	or (d287, d243, d251);
	xor (d288, d260, d277);
	or (d289, d251, d274);
	xor (d290, d243, d268);
	nor (d291, d243, d258);
	xnor (d292, d239, d263);
	nand (d293, d249, d251);
	or (d294, d250, d260);
	or (d295, d240, d252);
	assign f1 = d286;
	assign f2 = d284;
endmodule
