module CCGRCG90( x0, x1, x2, x3, f1, f2, f3, f4, f5, f6, f7, f8, f9 );

	input x0, x1, x2, x3;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109;

	buf (d1, x2);
	nor (d2, x0, x2);
	buf (d3, x1);
	not (d4, x0);
	not (d5, x2);
	or (d6, x2);
	nand (d7, x0);
	nand (d8, x1, x3);
	nand (d9, x0, x1);
	and (d10, x1, x2);
	and (d11, x1);
	xnor (d12, x3);
	nor (d13, x2);
	or (d14, x1);
	nor (d15, x1, x2);
	nor (d16, x0, x1);
	nor (d17, x2, x3);
	and (d18, x0);
	nand (d19, x3);
	xor (d20, x0, x3);
	or (d21, x1, x2);
	xnor (d22, x2, x3);
	or (d23, x2, x3);
	nand (d24, x0, x2);
	xnor (d25, x2);
	buf (d26, x0);
	xor (d27, x2);
	nor (d28, x0, x3);
	not (d29, x3);
	xnor (d30, x0);
	or (d31, x0, x2);
	xor (d32, x2, x3);
	xor (d33, x0, x1);
	or (d34, x0, x3);
	xnor (d35, x1);
	or (d36, x0, x1);
	or (d37, x1, x2);
	nor (d38, x0);
	nor (d39, x0, x3);
	xor (d40, x0);
	xor (d41, x1);
	and (d42, x2);
	nor (d43, x2, x3);
	not (d44, d39);
	nor (d45, d20, d30);
	nor (d46, d11, d17);
	nor (d47, d24, d39);
	nor (d48, d18, d25);
	buf (d49, d10);
	not (d50, d40);
	not (d51, d4);
	xnor (d52, d44, d45);
	xnor (d53, d46, d48);
	buf (d54, d23);
	nand (d55, d46, d48);
	nand (d56, d47, d48);
	nor (d57, d44, d45);
	xnor (d58, d46, d47);
	xor (d59, d44, d48);
	xnor (d60, d44);
	nor (d61, d44, d47);
	and (d62, d44, d46);
	not (d63, d14);
	nor (d64, d44, d48);
	nor (d65, d46, d48);
	or (d66, d44, d48);
	xor (d67, d47);
	and (d68, d45, d46);
	buf (d69, d30);
	buf (d70, d22);
	buf (d71, d36);
	nand (d72, d44, d46);
	and (d73, d48);
	xnor (d74, d44, d48);
	buf (d75, d32);
	xor (d76, d45, d47);
	not (d77, d47);
	nand (d78, d44);
	xnor (d79, d45, d48);
	and (d80, d45, d47);
	nor (d81, d46);
	buf (d82, d18);
	xnor (d83, d45, d47);
	or (d84, d46);
	nand (d85, d45, d48);
	nor (d86, d48);
	and (d87, d45, d48);
	xnor (d88, d45, d46);
	nand (d89, d47);
	nor (d90, d45, d47);
	and (d91, d45, d46);
	buf (d92, d31);
	nor (d93, d47, d48);
	xor (d94, d44, d48);
	nor (d95, d44, d48);
	nand (d96, d44, d46);
	buf (d97, d48);
	nor (d98, d45, d46);
	xnor (d99, d45, d48);
	and (d100, d46, d48);
	xor (d101, d45, d48);
	and (d102, d44, d47);
	xor (d103, d44, d45);
	buf (d104, d28);
	not (d105, d33);
	nand (d106, d45, d47);
	and (d107, d45, d48);
	buf (d108, d13);
	nor (d109, d44, d46);
	assign f1 = d104;
	assign f2 = d76;
	assign f3 = d64;
	assign f4 = d58;
	assign f5 = d81;
	assign f6 = d66;
	assign f7 = d108;
	assign f8 = d60;
	assign f9 = d76;
endmodule
