module CCGRCG114( x0, x1, x2, x3, x4, f1, f2 );

	input x0, x1, x2, x3, x4;
	output f1, f2;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133;

	nand (d1, x1, x2);
	nand (d2, x2, x3);
	and (d3, x2, x3);
	xnor (d4, x1, x4);
	nand (d5, x2, x4);
	buf (d6, x2);
	buf (d7, x4);
	not (d8, x2);
	xor (d9, x2, x3);
	nand (d10, d1);
	xor (d11, d4, d7);
	nor (d12, d2, d6);
	nor (d13, d4, d5);
	and (d14, d4, d7);
	not (d15, d9);
	nor (d16, d3, d7);
	buf (d17, d7);
	or (d18, d1, d3);
	nor (d19, d1, d6);
	buf (d20, d5);
	or (d21, d2);
	xnor (d22, d4, d5);
	xnor (d23, d2, d9);
	nand (d24, d2, d6);
	xnor (d25, d6, d7);
	nor (d26, d1, d5);
	and (d27, d2, d6);
	not (d28, d3);
	xnor (d29, d1, d4);
	nor (d30, d2, d3);
	or (d31, d4, d7);
	not (d32, d2);
	buf (d33, d9);
	buf (d34, x3);
	xor (d35, d5, d6);
	and (d36, d5, d8);
	xnor (d37, d2, d8);
	xnor (d38, d1, d7);
	xnor (d39, d1, d6);
	nor (d40, d1, d2);
	or (d41, d2, d4);
	or (d42, d22, d41);
	nor (d43, d30, d31);
	xor (d44, d28, d39);
	and (d45, d18, d39);
	xnor (d46, d12, d28);
	nand (d47, d14, d38);
	xor (d48, d15, d19);
	xor (d49, d14, d33);
	nor (d50, d20, d37);
	not (d51, d30);
	not (d52, d6);
	nand (d53, d26, d34);
	nor (d54, d32);
	xnor (d55, d14, d23);
	or (d56, d15, d33);
	or (d57, d19, d33);
	xnor (d58, d16, d38);
	xnor (d59, d22, d25);
	xor (d60, d19, d20);
	buf (d61, d15);
	buf (d62, d40);
	and (d63, d36, d38);
	nand (d64, d11, d25);
	xnor (d65, d17, d38);
	or (d66, d16, d22);
	nand (d67, d35, d37);
	and (d68, d20, d23);
	not (d69, d34);
	nor (d70, d24, d26);
	xor (d71, d12, d26);
	xnor (d72, d14, d19);
	buf (d73, d11);
	or (d74, d11, d13);
	nand (d75, d16, d21);
	not (d76, d40);
	and (d77, d11, d41);
	or (d78, d22, d36);
	nand (d79, d19, d30);
	and (d80, d14, d38);
	buf (d81, d21);
	and (d82, d12, d33);
	buf (d83, d26);
	or (d84, d16, d18);
	xnor (d85, d10, d31);
	and (d86, d22, d32);
	not (d87, d21);
	not (d88, d23);
	xor (d89, d26, d28);
	xor (d90, d16, d26);
	and (d91, d10, d41);
	and (d92, d12, d18);
	or (d93, d20, d36);
	nor (d94, d18, d32);
	nand (d95, d16, d38);
	buf (d96, d33);
	not (d97, x1);
	buf (d98, d17);
	buf (d99, d19);
	not (d100, d5);
	xnor (d101, d20, d40);
	xor (d102, d14, d24);
	nand (d103, d34, d36);
	buf (d104, d38);
	nand (d105, d35, d40);
	not (d106, d38);
	or (d107, d16, d21);
	buf (d108, d37);
	or (d109, d16, d28);
	nand (d110, d15, d36);
	and (d111, d36, d37);
	xor (d112, d24, d25);
	and (d113, d30, d41);
	xor (d114, d20, d25);
	not (d115, d14);
	xor (d116, d36, d39);
	nor (d117, d26, d39);
	buf (d118, d2);
	xor (d119, d19, d32);
	and (d120, d12, d29);
	not (d121, d31);
	and (d122, d26, d28);
	or (d123, d11, d27);
	and (d124, d25, d37);
	or (d125, d22, d38);
	buf (d126, d41);
	xor (d127, d14, d41);
	xor (d128, d33, d39);
	and (d129, d28, d38);
	not (d130, d26);
	and (d131, d25, d41);
	and (d132, d16, d27);
	not (d133, d32);
	assign f1 = d110;
	assign f2 = d81;
endmodule
