module CCGRCG113( x0, x1, x2, x3, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17, f18, f19, f20 );

	input x0, x1, x2, x3;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17, f18, f19, f20;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314, d315, d316, d317, d318, d319, d320, d321, d322, d323, d324, d325, d326, d327, d328, d329, d330, d331, d332, d333, d334, d335, d336, d337, d338, d339, d340, d341, d342, d343, d344, d345, d346, d347, d348, d349, d350, d351, d352, d353, d354, d355, d356, d357;

	nand (d1, x0, x1);
	nand (d2, x0, x2);
	nand (d3, x1);
	nand (d4, x1, x3);
	nand (d5, x2, x3);
	nand (d6, x1, x2);
	buf (d7, x2);
	or (d8, x0, x2);
	and (d9, x1, x3);
	xor (d10, x1);
	and (d11, x2, x3);
	xor (d12, x2, x3);
	xnor (d13, x0, x2);
	and (d14, x3);
	or (d15, x2, x3);
	xor (d16, d6, d14);
	nor (d17, d12, d15);
	buf (d18, x1);
	or (d19, d6, d14);
	not (d20, d11);
	or (d21, d6, d15);
	xnor (d22, d1, d7);
	and (d23, d9, d12);
	nor (d24, d2, d14);
	nor (d25, d8, d14);
	nor (d26, d3, d11);
	or (d27, d2, d15);
	buf (d28, d14);
	buf (d29, d13);
	buf (d30, d1);
	nor (d31, d5, d12);
	xnor (d32, d6, d15);
	xor (d33, d6, d11);
	and (d34, d9, d15);
	or (d35, d5, d10);
	nand (d36, d7, d14);
	nor (d37, d2, d14);
	xor (d38, d13, d15);
	or (d39, d12, d15);
	or (d40, d6, d11);
	buf (d41, d8);
	and (d42, d7, d13);
	nand (d43, d10, d14);
	not (d44, x2);
	xnor (d45, d11);
	nand (d46, d10, d14);
	buf (d47, d6);
	and (d48, d3, d15);
	not (d49, d5);
	xor (d50, d9, d15);
	nor (d51, d8, d15);
	and (d52, d9, d10);
	not (d53, d4);
	not (d54, d2);
	xor (d55, d7, d9);
	xor (d56, d2, d12);
	xnor (d57, d6, d8);
	xor (d58, d3, d6);
	nand (d59, d5, d14);
	xor (d60, d7, d10);
	nand (d61, d5, d6);
	not (d62, d7);
	nor (d63, d3, d13);
	and (d64, d2, d4);
	buf (d65, d3);
	not (d66, d10);
	nor (d67, d5, d13);
	buf (d68, d4);
	or (d69, d8, d11);
	xnor (d70, d6, d10);
	and (d71, d7, d10);
	and (d72, d3, d8);
	nand (d73, d2, d12);
	not (d74, x0);
	or (d75, d10);
	and (d76, d7, d12);
	nand (d77, d4, d12);
	not (d78, d6);
	or (d79, d42, d62);
	not (d80, d71);
	or (d81, d20, d51);
	xnor (d82, d38, d42);
	nor (d83, d30, d72);
	not (d84, d18);
	or (d85, d31, d63);
	nand (d86, d22, d62);
	and (d87, d29, d33);
	buf (d88, d56);
	buf (d89, d58);
	not (d90, d27);
	nand (d91, d55, d61);
	or (d92, d63, d74);
	xor (d93, d24, d55);
	xnor (d94, d38, d50);
	xor (d95, d33, d73);
	buf (d96, x3);
	and (d97, d29, d66);
	xnor (d98, d71, d73);
	nor (d99, d38, d48);
	xor (d100, d46, d50);
	xor (d101, d19, d72);
	not (d102, d16);
	or (d103, d48, d53);
	xor (d104, d64, d76);
	and (d105, d28, d65);
	nand (d106, d42, d62);
	nand (d107, d26, d56);
	or (d108, d20, d59);
	nor (d109, d45, d66);
	buf (d110, d30);
	nor (d111, d23, d52);
	or (d112, d18, d67);
	nand (d113, d22, d26);
	not (d114, d40);
	not (d115, d45);
	xnor (d116, d40, d68);
	nor (d117, d35, d73);
	xor (d118, d23, d51);
	nand (d119, d68, d73);
	or (d120, d58, d72);
	xnor (d121, d23, d46);
	xor (d122, d28, d54);
	xnor (d123, d34, d78);
	or (d124, d44, d66);
	nor (d125, d48, d69);
	nor (d126, d61, d65);
	not (d127, d28);
	not (d128, d78);
	nand (d129, d20, d42);
	or (d130, d43, d69);
	and (d131, d39, d76);
	and (d132, d46, d67);
	or (d133, d60, d66);
	xnor (d134, d59, d65);
	or (d135, d31, d72);
	nor (d136, d31, d70);
	xor (d137, d23, d33);
	nand (d138, d63);
	xnor (d139, d54, d59);
	xnor (d140, d67, d73);
	nand (d141, d29, d33);
	xor (d142, d34, d66);
	nor (d143, d22, d67);
	not (d144, d50);
	xnor (d145, d28, d74);
	xnor (d146, d62, d67);
	and (d147, d27, d34);
	buf (d148, d25);
	nand (d149, d54, d60);
	nand (d150, d35, d67);
	not (d151, d53);
	xnor (d152, d31, d40);
	or (d153, d33, d62);
	nand (d154, d34, d43);
	nor (d155, d59, d74);
	xor (d156, d32, d67);
	nor (d157, d67, d75);
	nand (d158, d31, d59);
	and (d159, d28, d57);
	nand (d160, d46, d53);
	buf (d161, d31);
	xnor (d162, d18, d20);
	nand (d163, d31, d39);
	nand (d164, d83, d109);
	and (d165, d107, d163);
	nand (d166, d101, d134);
	buf (d167, d131);
	and (d168, d80, d88);
	nor (d169, d110, d162);
	and (d170, d90, d93);
	and (d171, d95, d122);
	xnor (d172, d103, d104);
	not (d173, d135);
	xor (d174, d79, d126);
	xnor (d175, d131, d161);
	xnor (d176, d89, d113);
	or (d177, d138, d158);
	xor (d178, d94, d136);
	nand (d179, d80, d85);
	nor (d180, d133, d155);
	nor (d181, d83, d128);
	buf (d182, d138);
	buf (d183, d152);
	buf (d184, d87);
	not (d185, d123);
	xor (d186, d83, d156);
	and (d187, d169, d183);
	xnor (d188, d165, d180);
	not (d189, d148);
	nor (d190, d169, d184);
	buf (d191, d167);
	or (d192, d171, d179);
	nand (d193, d166, d183);
	xnor (d194, d169, d178);
	not (d195, d22);
	xnor (d196, d165, d175);
	or (d197, d172, d183);
	nand (d198, d174, d178);
	and (d199, d182, d183);
	xnor (d200, d167, d177);
	xor (d201, d167, d179);
	or (d202, d165, d171);
	nor (d203, d165, d177);
	xor (d204, d172, d185);
	or (d205, d172, d180);
	xor (d206, d173, d184);
	not (d207, d49);
	xor (d208, d178, d179);
	or (d209, d172, d181);
	not (d210, d153);
	xnor (d211, d166, d169);
	buf (d212, d83);
	xnor (d213, d178, d180);
	nand (d214, d164, d168);
	nor (d215, d170, d185);
	and (d216, d171, d183);
	nor (d217, d181, d183);
	and (d218, d170, d172);
	xor (d219, d168, d176);
	nor (d220, d166, d182);
	buf (d221, d62);
	nand (d222, d172, d183);
	or (d223, d201, d207);
	and (d224, d189, d207);
	xnor (d225, d192, d218);
	or (d226, d190, d191);
	xnor (d227, d201, d205);
	xor (d228, d195, d201);
	nor (d229, d190, d192);
	nand (d230, d200, d208);
	xor (d231, d199, d214);
	xor (d232, d194, d217);
	xor (d233, d196, d215);
	xnor (d234, d187, d196);
	or (d235, d197, d208);
	or (d236, d200, d219);
	xor (d237, d200);
	xnor (d238, d210, d214);
	or (d239, d215, d216);
	nand (d240, d191, d192);
	nand (d241, d215, d221);
	nand (d242, d206, d222);
	nand (d243, d193, d196);
	nor (d244, d206, d212);
	xor (d245, d198, d207);
	not (d246, d93);
	xnor (d247, d212, d222);
	not (d248, d80);
	not (d249, d70);
	and (d250, d190, d214);
	or (d251, d195, d196);
	xnor (d252, d188, d203);
	nand (d253, d191, d211);
	or (d254, d212, d218);
	nand (d255, d188, d206);
	or (d256, d206, d212);
	xor (d257, d206, d220);
	or (d258, d200, d204);
	buf (d259, d100);
	xor (d260, d199, d219);
	nor (d261, d208, d209);
	xnor (d262, d187, d210);
	and (d263, d194, d201);
	nor (d264, d212, d219);
	buf (d265, d124);
	nor (d266, d194, d205);
	or (d267, d200, d222);
	not (d268, d81);
	not (d269, d103);
	not (d270, d216);
	xnor (d271, d200, d213);
	not (d272, d12);
	xor (d273, d203, d213);
	nand (d274, d190, d211);
	buf (d275, d75);
	nand (d276, d207, d220);
	and (d277, d207, d216);
	and (d278, d208, d210);
	nor (d279, d188, d217);
	and (d280, d197, d216);
	nand (d281, d190, d207);
	nor (d282, d197, d206);
	buf (d283, d96);
	xnor (d284, d199, d220);
	and (d285, d188, d212);
	nor (d286, d200, d222);
	or (d287, d193, d197);
	nand (d288, d188, d218);
	nand (d289, d187, d200);
	or (d290, d192, d208);
	nand (d291, d270, d278);
	and (d292, d231);
	buf (d293, d97);
	xor (d294, d242, d251);
	not (d295, d193);
	nand (d296, d266, d271);
	nor (d297, d224, d255);
	nand (d298, d228, d247);
	or (d299, d245, d286);
	or (d300, d230, d266);
	nor (d301, d250, d252);
	or (d302, d225, d287);
	not (d303, d94);
	buf (d304, d285);
	xnor (d305, d255, d290);
	and (d306, d228, d231);
	nor (d307, d240, d256);
	or (d308, d228, d249);
	xor (d309, d280, d281);
	xnor (d310, d224, d225);
	xnor (d311, d259, d266);
	xnor (d312, d225, d261);
	xnor (d313, d229, d240);
	nor (d314, d242, d257);
	buf (d315, d92);
	and (d316, d302, d314);
	and (d317, d299, d309);
	not (d318, d41);
	or (d319, d309, d314);
	nor (d320, d309, d314);
	or (d321, d291, d296);
	nand (d322, d300, d308);
	and (d323, d292, d297);
	buf (d324, d259);
	and (d325, d291, d315);
	or (d326, d295, d315);
	nor (d327, d302);
	or (d328, d297, d305);
	nor (d329, d292, d309);
	xnor (d330, d291, d312);
	not (d331, d87);
	not (d332, d152);
	not (d333, d298);
	xor (d334, d295, d296);
	xor (d335, d297, d311);
	nand (d336, d308, d315);
	and (d337, d292, d308);
	nor (d338, d300, d302);
	xnor (d339, d292, d300);
	nand (d340, d295, d302);
	nor (d341, d293, d304);
	and (d342, d307, d315);
	xnor (d343, d300, d301);
	and (d344, d301, d306);
	xnor (d345, d307, d308);
	and (d346, d291, d305);
	not (d347, d74);
	nand (d348, d297, d299);
	nand (d349, d295, d314);
	or (d350, d295, d296);
	not (d351, d194);
	not (d352, d157);
	or (d353, d305, d313);
	buf (d354, d239);
	not (d355, d26);
	or (d356, d300, d307);
	xnor (d357, d294, d309);
	assign f1 = d348;
	assign f2 = d321;
	assign f3 = d340;
	assign f4 = d342;
	assign f5 = d324;
	assign f6 = d334;
	assign f7 = d316;
	assign f8 = d319;
	assign f9 = d321;
	assign f10 = d316;
	assign f11 = d337;
	assign f12 = d331;
	assign f13 = d353;
	assign f14 = d351;
	assign f15 = d343;
	assign f16 = d345;
	assign f17 = d342;
	assign f18 = d317;
	assign f19 = d343;
	assign f20 = d354;
endmodule
