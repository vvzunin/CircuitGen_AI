module CCGRCG189( x0, x1, x2, x3, x4, x5, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17, f18, f19, f20 );

	input x0, x1, x2, x3, x4, x5;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17, f18, f19, f20;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240;

	nor (d1, x3, x5);
	and (d2, x1, x3);
	buf (d3, x2);
	or (d4, x2, x3);
	nand (d5, x2, x5);
	and (d6, x1, x2);
	xor (d7, x0, x1);
	xnor (d8, x3, x5);
	or (d9, x0, x4);
	xnor (d10, x2, x5);
	or (d11, x1, x5);
	not (d12, x3);
	buf (d13, x1);
	xor (d14, x1);
	xor (d15, x2, x3);
	xnor (d16, x0, x1);
	or (d17, x1, x5);
	xor (d18, x3, x5);
	and (d19, x0, x1);
	nand (d20, x5);
	not (d21, x1);
	xnor (d22, x1, x2);
	xnor (d23, x2, x5);
	xnor (d24, x3);
	xnor (d25, x4, x5);
	and (d26, x4);
	nand (d27, x4);
	xor (d28, x2, x4);
	nor (d29, x4, x5);
	nor (d30, x2, x3);
	nor (d31, x0, x1);
	and (d32, x1, x3);
	xor (d33, x0, x1);
	and (d34, x2, x4);
	and (d35, x3, x5);
	not (d36, x4);
	nand (d37, x0);
	or (d38, x0, x3);
	not (d39, x2);
	or (d40, x0);
	xor (d41, x1, x2);
	xnor (d42, x1);
	not (d43, x0);
	nand (d44, x3, x4);
	nand (d45, x2, x5);
	and (d46, x3);
	or (d47, x1, x3);
	and (d48, x3, x5);
	and (d49, x2);
	nor (d50, x3, x5);
	nand (d51, x0, x2);
	xor (d52, x3, x5);
	or (d53, x2, x4);
	or (d54, x3, x4);
	and (d55, x0, x3);
	xor (d56, x0, x4);
	and (d57, x1, x5);
	xnor (d58, x0, x2);
	xnor (d59, x0, x5);
	buf (d60, x3);
	xor (d61, x3, x4);
	xnor (d62, d46, d59);
	xor (d63, d35, d59);
	buf (d64, d15);
	and (d65, d38, d61);
	nand (d66, d25, d58);
	xor (d67, d3, d21);
	xnor (d68, d20, d23);
	not (d69, d22);
	nor (d70, d1, d14);
	xnor (d71, d10);
	not (d72, d53);
	xor (d73, d14, d28);
	nor (d74, d19, d20);
	xor (d75, d22, d25);
	xor (d76, d40, d54);
	not (d77, d7);
	xnor (d78, d1, d41);
	buf (d79, d57);
	nand (d80, d36, d48);
	nor (d81, d65, d75);
	xnor (d82, d62, d72);
	buf (d83, d73);
	xor (d84, d78, d80);
	xnor (d85, d71, d78);
	buf (d86, d55);
	not (d87, d35);
	not (d88, d75);
	buf (d89, d74);
	nor (d90, d65, d77);
	not (d91, d79);
	and (d92, d64, d72);
	xor (d93, d71, d72);
	or (d94, d62, d74);
	xnor (d95, d67, d78);
	not (d96, d11);
	not (d97, d56);
	and (d98, d62, d68);
	and (d99, d69, d78);
	xnor (d100, d62, d66);
	nor (d101, d69, d70);
	nand (d102, d72, d78);
	or (d103, d67, d73);
	and (d104, d63, d67);
	buf (d105, d33);
	and (d106, d76, d77);
	nand (d107, d75, d77);
	buf (d108, d35);
	not (d109, d45);
	and (d110, d63, d75);
	not (d111, d50);
	and (d112, d69, d75);
	and (d113, d72, d80);
	nor (d114, d68, d76);
	nor (d115, d76, d79);
	nor (d116, d67, d73);
	nand (d117, d64, d76);
	xor (d118, d63, d66);
	or (d119, d62, d75);
	and (d120, d66, d73);
	or (d121, d71, d72);
	nand (d122, d63, d78);
	nor (d123, d78, d80);
	nand (d124, d62, d76);
	buf (d125, d49);
	and (d126, d64, d75);
	xnor (d127, d74, d77);
	and (d128, d70, d73);
	nor (d129, d64, d78);
	and (d130, d68, d69);
	nor (d131, d64, d65);
	xor (d132, d79, d80);
	nor (d133, d76, d78);
	not (d134, d12);
	not (d135, d54);
	nor (d136, d69, d75);
	xor (d137, d74);
	nor (d138, d64, d71);
	not (d139, d61);
	xor (d140, d67, d77);
	and (d141, d74, d76);
	and (d142, d73, d78);
	xnor (d143, d66, d67);
	nand (d144, d63, d74);
	xor (d145, d65, d73);
	xor (d146, d62, d73);
	xnor (d147, d67, d75);
	not (d148, d4);
	or (d149, d68, d75);
	nand (d150, d67, d72);
	nand (d151, d69, d78);
	or (d152, d77, d80);
	buf (d153, d2);
	xnor (d154, d65, d66);
	and (d155, d64, d69);
	nand (d156, d71, d80);
	buf (d157, d25);
	nor (d158, d66, d76);
	and (d159, d97, d156);
	buf (d160, d27);
	or (d161, d115, d149);
	not (d162, d154);
	nand (d163, d134, d138);
	and (d164, d83, d114);
	xor (d165, d96, d122);
	xnor (d166, d114, d156);
	not (d167, d98);
	not (d168, d109);
	nand (d169, d82, d96);
	and (d170, d98, d149);
	buf (d171, d134);
	xor (d172, d81, d84);
	nor (d173, d149, d150);
	buf (d174, d69);
	buf (d175, d149);
	nand (d176, d88, d95);
	xnor (d177, d85, d110);
	nand (d178, d111, d155);
	nand (d179, d105, d114);
	not (d180, d158);
	or (d181, d111, d140);
	xor (d182, d82, d125);
	nor (d183, d110, d156);
	and (d184, d123, d156);
	buf (d185, d119);
	buf (d186, d58);
	xnor (d187, d95, d113);
	and (d188, d87, d146);
	not (d189, d143);
	not (d190, d48);
	or (d191, d145);
	xor (d192, d98, d109);
	xor (d193, d119, d134);
	not (d194, d34);
	xor (d195, d114, d157);
	xor (d196, d105, d144);
	nor (d197, d108, d141);
	xnor (d198, d149, d155);
	or (d199, d118, d129);
	or (d200, d132, d151);
	not (d201, d78);
	not (d202, d130);
	and (d203, d102, d107);
	or (d204, d90, d99);
	nand (d205, d84, d145);
	not (d206, d119);
	xnor (d207, d92, d102);
	buf (d208, d54);
	or (d209, d96, d144);
	nor (d210, d96, d121);
	xnor (d211, d165, d197);
	nand (d212, d173, d204);
	and (d213, d189, d192);
	not (d214, d51);
	nor (d215, d198, d208);
	not (d216, d95);
	or (d217, d165, d166);
	and (d218, d216, d217);
	xor (d219, d213);
	buf (d220, d70);
	xnor (d221, d211, d212);
	or (d222, d211, d212);
	not (d223, d24);
	and (d224, d213, d215);
	nand (d225, d214, d217);
	nand (d226, d212, d215);
	nand (d227, d214, d217);
	nor (d228, d216, d217);
	xnor (d229, d213, d214);
	xor (d230, d212, d216);
	buf (d231, d194);
	nor (d232, d211, d215);
	buf (d233, d68);
	not (d234, d125);
	nand (d235, d212, d217);
	xor (d236, d211, d213);
	buf (d237, d92);
	or (d238, d213, d216);
	xor (d239, d211, d212);
	xor (d240, d212);
	assign f1 = d237;
	assign f2 = d224;
	assign f3 = d219;
	assign f4 = d237;
	assign f5 = d229;
	assign f6 = d240;
	assign f7 = d231;
	assign f8 = d237;
	assign f9 = d219;
	assign f10 = d227;
	assign f11 = d230;
	assign f12 = d218;
	assign f13 = d225;
	assign f14 = d238;
	assign f15 = d219;
	assign f16 = d223;
	assign f17 = d226;
	assign f18 = d222;
	assign f19 = d233;
	assign f20 = d224;
endmodule
