// Benchmark "CCGRCG165" written by ABC on Tue Feb 13 20:52:15 2024

module CCGRCG165 ( 
    x0, x1, x2, x3, x4, x5,
    f1, f2, f3, f4, f5, f6, f7, f8  );
  input  x0, x1, x2, x3, x4, x5;
  output f1, f2, f3, f4, f5, f6, f7, f8;
  wire new_n15_, new_n16_, new_n18_, new_n20_, new_n23_, new_n24_;
  assign new_n15_ = ~x0 & ~x1;
  assign new_n16_ = x0 & x1;
  assign f1 = ~new_n15_ & ~new_n16_;
  assign new_n18_ = x0 & x4;
  assign f2 = ~new_n18_;
  assign new_n20_ = ~x0 & ~x4;
  assign f3 = ~new_n20_ & ~new_n18_;
  assign f4 = x0 & x5;
  assign new_n23_ = ~x3 & ~x5;
  assign new_n24_ = x3 & x5;
  assign f6 = ~new_n23_ & ~new_n24_;
  assign f8 = ~x2 & ~x5;
  assign f5 = x5;
  assign f7 = x0;
endmodule


