module CCGRCG3( x0, x1, f1, f2 );

	input x0, x1;
	output f1, f2;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147;

	xnor (d1, x0, x1);
	xor (d2, x1);
	nor (d3, x0, x1);
	not (d4, x1);
	buf (d5, x0);
	nor (d6, x0, x1);
	and (d7, x1);
	and (d8, x0, x1);
	xor (d9, x0, x1);
	or (d10, x0);
	nand (d11, x0, x1);
	buf (d12, x1);
	or (d13, x0, x1);
	or (d14, x1);
	xor (d15, x0);
	nand (d16, x1);
	or (d17, x0, x1);
	xnor (d18, x0, x1);
	xnor (d19, x1);
	and (d20, x0, x1);
	xor (d21, x0, x1);
	nand (d22, x0);
	nand (d23, x0, x1);
	xnor (d24, x0);
	and (d25, x0);
	nor (d26, x0);
	and (d27, d13, d23);
	nor (d28, d6, d23);
	buf (d29, d10);
	xnor (d30, d9, d13);
	or (d31, d7, d21);
	nand (d32, d12, d21);
	xor (d33, d1, d16);
	xnor (d34, d2, d11);
	and (d35, d11, d19);
	nand (d36, d10, d11);
	xor (d37, d1, d3);
	xor (d38, d7, d16);
	not (d39, d4);
	nor (d40, d4, d19);
	xnor (d41, d12, d14);
	or (d42, d12, d18);
	or (d43, d14, d19);
	buf (d44, d1);
	xnor (d45, d10, d11);
	or (d46, d3, d24);
	and (d47, d10, d15);
	nor (d48, d10, d24);
	buf (d49, d12);
	xnor (d50, d3, d16);
	not (d51, d1);
	not (d52, d3);
	nand (d53, d9, d20);
	nand (d54, d13, d22);
	and (d55, d11, d23);
	buf (d56, d13);
	not (d57, d11);
	nor (d58, d1, d3);
	xor (d59, d1, d19);
	nand (d60, d27, d43);
	buf (d61, d18);
	not (d62, d32);
	xor (d63, d42, d44);
	not (d64, d23);
	or (d65, d46, d49);
	nand (d66, d27, d46);
	and (d67, d40, d51);
	nor (d68, d45, d57);
	and (d69, d45, d59);
	or (d70, d27, d45);
	xor (d71, d31, d58);
	xnor (d72, d36, d58);
	nand (d73, d40, d44);
	not (d74, d8);
	nand (d75, d33, d45);
	xor (d76, d27, d35);
	and (d77, d42);
	nor (d78, d31, d40);
	xor (d79, d48, d51);
	nor (d80, d33, d52);
	nand (d81, d35, d42);
	or (d82, d36, d59);
	buf (d83, d5);
	buf (d84, d40);
	xor (d85, d36, d39);
	xnor (d86, d30, d47);
	buf (d87, d9);
	xor (d88, d39, d56);
	not (d89, d18);
	or (d90, d50, d56);
	xnor (d91, d27, d46);
	nand (d92, d41, d42);
	and (d93, d48, d50);
	and (d94, d52, d56);
	nand (d95, d38, d47);
	or (d96, d39, d43);
	xnor (d97, d37, d38);
	nor (d98, d30, d52);
	or (d99, d29, d58);
	or (d100, d42, d52);
	buf (d101, d20);
	or (d102, d40, d44);
	nand (d103, d30, d59);
	xnor (d104, d29);
	xor (d105, d56, d58);
	buf (d106, d65);
	and (d107, d60, d64);
	xor (d108, d78, d99);
	or (d109, d64, d103);
	buf (d110, d78);
	nor (d111, d79, d102);
	not (d112, d62);
	xnor (d113, d61, d98);
	and (d114, d62, d99);
	and (d115, d90, d102);
	buf (d116, d30);
	nor (d117, d85, d102);
	xor (d118, d72, d75);
	nor (d119, d68, d72);
	nor (d120, d76, d100);
	xor (d121, d101, d105);
	and (d122, d78, d87);
	not (d123, d36);
	xnor (d124, d77, d101);
	buf (d125, d59);
	nor (d126, d61, d96);
	xnor (d127, d67, d74);
	buf (d128, d67);
	and (d129, d78, d81);
	xnor (d130, d60, d105);
	or (d131, d72, d105);
	nor (d132, d92, d105);
	and (d133, d101, d105);
	buf (d134, d73);
	not (d135, d81);
	nand (d136, d77, d92);
	xnor (d137, d62, d95);
	nand (d138, d60, d99);
	buf (d139, d34);
	or (d140, d63, d69);
	not (d141, d86);
	or (d142, d67, d70);
	xnor (d143, d63, d93);
	or (d144, d75, d99);
	or (d145, d60, d61);
	xor (d146, d82, d100);
	not (d147, d51);
	assign f1 = d111;
	assign f2 = d110;
endmodule
