module CCGRCG161( x0, x1, x2, x3, x4, x5, f1, f2, f3, f4, f5, f6 );

	input x0, x1, x2, x3, x4, x5;
	output f1, f2, f3, f4, f5, f6;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314, d315, d316, d317, d318, d319, d320, d321, d322, d323, d324, d325, d326, d327, d328, d329, d330, d331, d332, d333, d334, d335, d336, d337, d338, d339, d340, d341, d342, d343, d344, d345, d346, d347, d348, d349, d350, d351, d352, d353, d354, d355, d356, d357, d358, d359, d360, d361, d362, d363, d364, d365, d366, d367, d368, d369, d370, d371, d372, d373, d374, d375, d376, d377, d378, d379, d380, d381, d382, d383, d384, d385, d386, d387, d388, d389, d390, d391, d392, d393, d394, d395, d396, d397, d398, d399, d400, d401, d402, d403, d404, d405, d406, d407, d408, d409, d410, d411, d412, d413, d414, d415, d416, d417, d418, d419, d420, d421, d422, d423, d424, d425, d426, d427, d428, d429, d430, d431, d432, d433, d434, d435, d436, d437, d438, d439, d440, d441, d442, d443, d444, d445;

	buf (d1, x1);
	xor (d2, x2, x3);
	buf (d3, x2);
	xnor (d4, x2, x4);
	and (d5, x0, x5);
	buf (d6, x4);
	xnor (d7, x1, x4);
	xor (d8, x0, x2);
	or (d9, x1, x4);
	not (d10, x1);
	nor (d11, x0);
	xor (d12, x1, x2);
	or (d13, x0);
	nand (d14, x2, x3);
	and (d15, x2, x4);
	nand (d16, x1, x4);
	not (d17, x3);
	buf (d18, x3);
	nor (d19, x1, x2);
	nor (d20, x3, x4);
	xor (d21, x0, x4);
	xnor (d22, x0);
	nor (d23, x0, x3);
	xnor (d24, x2, x5);
	and (d25, x1);
	xor (d26, x2, x4);
	xor (d27, x0, x1);
	xor (d28, x1, x5);
	and (d29, x1, x2);
	and (d30, x2, x5);
	nor (d31, x0, x2);
	nand (d32, x0, x5);
	and (d33, x4);
	or (d34, x4);
	xnor (d35, x1, x3);
	or (d36, x0, x4);
	xnor (d37, x4, x5);
	nor (d38, x0, x4);
	xnor (d39, x2, x5);
	xor (d40, x0, x5);
	nor (d41, x3, x4);
	nor (d42, x1, x3);
	and (d43, x2, x3);
	nand (d44, x0, x4);
	not (d45, x4);
	nor (d46, x2, x4);
	xor (d47, x0, x3);
	or (d48, x1, x5);
	xnor (d49, x2, x4);
	nand (d50, x0, x3);
	xnor (d51, x3, x5);
	buf (d52, x0);
	nand (d53, x0, x1);
	and (d54, x5);
	and (d55, x0, x1);
	xnor (d56, x1, x2);
	not (d57, x5);
	buf (d58, x5);
	nor (d59, x0, x3);
	nand (d60, x0, x2);
	nand (d61, x2, x4);
	and (d62, x3, x5);
	xnor (d63, x3, x5);
	nand (d64, x0);
	nand (d65, x0, x5);
	or (d66, x2);
	nand (d67, x1, x5);
	xor (d68, d12, d28);
	and (d69, d46, d52);
	or (d70, d45, d60);
	buf (d71, d20);
	or (d72, d46, d48);
	and (d73, d25, d38);
	and (d74, d2, d7);
	and (d75, d28, d62);
	nor (d76, d28, d40);
	xor (d77, d38, d47);
	or (d78, d21, d30);
	xnor (d79, d69, d72);
	nor (d80, d70, d71);
	nand (d81, d68, d72);
	nor (d82, d72, d73);
	buf (d83, d45);
	xor (d84, d69, d70);
	not (d85, d65);
	xnor (d86, d75);
	xor (d87, d70, d77);
	buf (d88, d32);
	nor (d89, d72, d74);
	xor (d90, d68, d76);
	nor (d91, d75, d77);
	not (d92, d49);
	nor (d93, d76, d77);
	xor (d94, d68, d69);
	nor (d95, d68, d74);
	xnor (d96, d70, d76);
	nand (d97, d68, d71);
	buf (d98, d1);
	buf (d99, d74);
	or (d100, d69, d74);
	not (d101, d53);
	not (d102, d33);
	buf (d103, d10);
	or (d104, d71);
	xnor (d105, d70, d72);
	nor (d106, d74, d78);
	or (d107, d73, d76);
	buf (d108, d56);
	nand (d109, d102, d104);
	and (d110, d102, d106);
	xnor (d111, d92, d93);
	xor (d112, d82, d85);
	xor (d113, d85, d89);
	or (d114, d83, d100);
	xor (d115, d86, d93);
	not (d116, d22);
	nand (d117, d92, d94);
	nand (d118, d86, d87);
	or (d119, d80, d100);
	buf (d120, d98);
	and (d121, d83, d87);
	not (d122, d86);
	nor (d123, d80, d105);
	buf (d124, d71);
	xor (d125, d79, d99);
	and (d126, d89, d101);
	buf (d127, d33);
	xor (d128, d84, d98);
	not (d129, d50);
	buf (d130, d31);
	xor (d131, d86, d102);
	buf (d132, d96);
	xnor (d133, d81, d87);
	nor (d134, d85, d95);
	xnor (d135, d83, d96);
	xor (d136, d85, d86);
	and (d137, d82, d95);
	xor (d138, d81, d95);
	nand (d139, d80, d85);
	nor (d140, d93, d101);
	xnor (d141, d83, d92);
	or (d142, d79, d88);
	not (d143, d15);
	xnor (d144, d90, d95);
	nand (d145, d79);
	nor (d146, d90, d94);
	or (d147, d85, d104);
	nand (d148, d91, d94);
	not (d149, d91);
	or (d150, d100, d107);
	buf (d151, d51);
	nand (d152, d86, d99);
	buf (d153, d25);
	nand (d154, d82, d87);
	nor (d155, d86, d98);
	or (d156, d91, d104);
	buf (d157, d107);
	or (d158, d79, d86);
	xnor (d159, d81, d92);
	and (d160, d89, d98);
	and (d161, d82, d106);
	nand (d162, d88, d95);
	xnor (d163, d82, d103);
	nand (d164, d86, d90);
	or (d165, d84, d93);
	or (d166, d103, d105);
	or (d167, d81, d86);
	nor (d168, d79);
	buf (d169, d2);
	buf (d170, d14);
	nand (d171, d100, d107);
	xor (d172, d102, d105);
	xor (d173, d80, d86);
	xnor (d174, d87, d106);
	xor (d175, d89, d106);
	xnor (d176, d91, d92);
	or (d177, d90, d92);
	xnor (d178, d91, d100);
	not (d179, d19);
	or (d180, d99, d101);
	and (d181, d85, d95);
	xnor (d182, d82);
	or (d183, d87);
	nor (d184, d91, d95);
	xor (d185, d94, d95);
	xor (d186, d79, d96);
	or (d187, d81, d92);
	not (d188, d36);
	not (d189, d67);
	xor (d190, d97, d103);
	buf (d191, d47);
	xor (d192, d134, d186);
	xnor (d193, d123, d157);
	nand (d194, d114, d146);
	buf (d195, d84);
	xnor (d196, d147, d163);
	xor (d197, d138, d161);
	not (d198, d48);
	nand (d199, d116, d181);
	xor (d200, d162, d187);
	not (d201, d173);
	nand (d202, d121, d172);
	buf (d203, d114);
	and (d204, d166, d173);
	xnor (d205, d111, d169);
	nand (d206, d146, d166);
	buf (d207, d183);
	xor (d208, d113, d176);
	nor (d209, d129, d164);
	xnor (d210, d134, d176);
	nor (d211, d119, d149);
	buf (d212, d61);
	or (d213, d147, d178);
	or (d214, d145, d191);
	nor (d215, d127, d161);
	nand (d216, d118, d165);
	nand (d217, d115, d165);
	nor (d218, d130, d150);
	nor (d219, d143, d160);
	nand (d220, d207, d215);
	nor (d221, d202, d217);
	nor (d222, d194, d202);
	nand (d223, d211, d215);
	and (d224, d200, d212);
	or (d225, d205, d219);
	nor (d226, d195, d216);
	not (d227, d169);
	or (d228, d206, d212);
	xor (d229, d193, d215);
	or (d230, d211, d215);
	buf (d231, d213);
	xnor (d232, d198, d213);
	nor (d233, d195, d212);
	not (d234, d141);
	nand (d235, d194, d203);
	xnor (d236, d194, d202);
	or (d237, d195, d205);
	xnor (d238, d207, d219);
	nand (d239, d192, d207);
	nand (d240, d203, d219);
	xor (d241, d210, d212);
	buf (d242, d205);
	nor (d243, d212, d219);
	and (d244, d206, d207);
	xor (d245, d209, d218);
	xor (d246, d202, d204);
	nor (d247, d193, d211);
	or (d248, d225, d241);
	xnor (d249, d233, d234);
	nor (d250, d227, d230);
	and (d251, d221, d229);
	nor (d252, d221, d224);
	buf (d253, d198);
	and (d254, d220, d233);
	nor (d255, d224, d239);
	nand (d256, d224, d230);
	xor (d257, d233, d239);
	xnor (d258, d242, d243);
	buf (d259, d69);
	nand (d260, d228, d247);
	xnor (d261, d232, d233);
	or (d262, d227, d230);
	buf (d263, d22);
	nor (d264, d238, d247);
	nand (d265, d222, d242);
	nor (d266, d222, d245);
	nand (d267, d220, d234);
	xor (d268, d222, d232);
	nor (d269, d241, d245);
	buf (d270, d75);
	xor (d271, d223, d226);
	xor (d272, d231, d239);
	not (d273, d183);
	nand (d274, d227, d246);
	nand (d275, d234, d243);
	or (d276, d235);
	or (d277, d237, d247);
	xor (d278, d228, d239);
	not (d279, d138);
	buf (d280, d200);
	and (d281, d229, d236);
	or (d282, d230, d245);
	and (d283, d229, d246);
	xor (d284, d233, d234);
	nor (d285, d251, d265);
	and (d286, d249, d251);
	nand (d287, d267, d279);
	nor (d288, d254, d282);
	nand (d289, d258, d283);
	xor (d290, d256, d266);
	buf (d291, d195);
	nand (d292, d270, d281);
	buf (d293, d41);
	nand (d294, d248, d260);
	xor (d295, d259, d270);
	or (d296, d248, d284);
	and (d297, d275, d278);
	or (d298, d249, d277);
	nand (d299, d271, d277);
	or (d300, d254, d284);
	xor (d301, d259, d275);
	not (d302, d51);
	xor (d303, d264, d279);
	and (d304, d253, d262);
	nor (d305, d254, d270);
	nand (d306, d273, d282);
	and (d307, d264, d274);
	or (d308, d269, d284);
	and (d309, d254, d278);
	xor (d310, d281, d283);
	xnor (d311, d266, d279);
	xor (d312, d270, d273);
	xor (d313, d251, d281);
	buf (d314, d260);
	nand (d315, d254, d255);
	not (d316, d18);
	and (d317, d251, d254);
	and (d318, d267, d270);
	nand (d319, d258, d275);
	xor (d320, d259, d262);
	nor (d321, d266, d269);
	nor (d322, d255, d274);
	nor (d323, d272, d274);
	nor (d324, d253, d259);
	and (d325, d254);
	nor (d326, d258, d265);
	or (d327, d258, d278);
	not (d328, d267);
	xor (d329, d281);
	or (d330, d267, d276);
	buf (d331, d143);
	not (d332, d299);
	xor (d333, d300, d304);
	xnor (d334, d287, d290);
	xnor (d335, d302, d325);
	xor (d336, d289, d312);
	xor (d337, d303, d321);
	nand (d338, d305, d315);
	xnor (d339, d304, d317);
	nand (d340, d298, d308);
	not (d341, d82);
	buf (d342, d315);
	or (d343, d308, d319);
	xor (d344, d305, d314);
	not (d345, d216);
	xnor (d346, d320, d322);
	not (d347, d205);
	or (d348, d310, d319);
	or (d349, d300, d328);
	xor (d350, d310, d324);
	or (d351, d322, d325);
	xnor (d352, d296, d302);
	xnor (d353, d287, d323);
	nand (d354, d291, d317);
	xnor (d355, d310, d315);
	xor (d356, d312, d313);
	xor (d357, d316, d319);
	nor (d358, d295, d306);
	or (d359, d296, d328);
	nor (d360, d317);
	not (d361, d68);
	and (d362, d302, d326);
	or (d363, d298, d319);
	nor (d364, d298, d324);
	not (d365, d130);
	not (d366, d111);
	and (d367, d310, d322);
	buf (d368, d37);
	buf (d369, d312);
	and (d370, d295, d329);
	or (d371, d285, d300);
	or (d372, d308, d317);
	nand (d373, d302, d312);
	or (d374, d292, d324);
	and (d375, d296, d330);
	xnor (d376, d294, d295);
	not (d377, d324);
	buf (d378, d29);
	not (d379, d285);
	nand (d380, d294, d325);
	or (d381, d293, d294);
	xnor (d382, d308, d320);
	buf (d383, d229);
	xor (d384, d286, d331);
	or (d385, d326, d330);
	nand (d386, d308, d330);
	nand (d387, d302, d303);
	nand (d388, d305, d321);
	nor (d389, d303, d317);
	xor (d390, d285, d323);
	nor (d391, d311, d330);
	buf (d392, d239);
	not (d393, d146);
	nor (d394, d307, d325);
	nor (d395, d294, d329);
	xnor (d396, d324, d325);
	and (d397, d313, d330);
	not (d398, d76);
	xnor (d399, d316, d331);
	nand (d400, d296, d326);
	buf (d401, d217);
	buf (d402, d97);
	and (d403, d292, d321);
	nand (d404, d327, d328);
	nor (d405, d301, d323);
	buf (d406, d154);
	or (d407, d335, d351);
	xor (d408, d355, d361);
	nor (d409, d354, d361);
	not (d410, d284);
	nor (d411, d360, d393);
	nand (d412, d343, d371);
	xnor (d413, d332, d346);
	nand (d414, d341, d364);
	not (d415, d165);
	and (d416, d332, d339);
	nand (d417, d392, d401);
	and (d418, d357, d365);
	xnor (d419, d388, d399);
	nor (d420, d371, d396);
	and (d421, d348, d403);
	nand (d422, d383, d388);
	nor (d423, d336, d347);
	and (d424, d335, d383);
	buf (d425, d216);
	nor (d426, d338, d357);
	xnor (d427, d366, d376);
	or (d428, d368, d385);
	not (d429, d393);
	not (d430, d309);
	nor (d431, d352, d392);
	nor (d432, d366, d375);
	nor (d433, d381, d382);
	or (d434, d355, d399);
	not (d435, d56);
	buf (d436, d332);
	nand (d437, d336, d395);
	xnor (d438, d388, d404);
	and (d439, d355, d385);
	or (d440, d358, d389);
	not (d441, d135);
	nand (d442, d398);
	or (d443, d358, d402);
	xor (d444, d364, d366);
	nand (d445, d363);
	assign f1 = d408;
	assign f2 = d417;
	assign f3 = d407;
	assign f4 = d441;
	assign f5 = d440;
	assign f6 = d427;
endmodule
