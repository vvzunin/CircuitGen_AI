module CCGRCG43( x0, x1, x2, x3, f1, f2 );

	input x0, x1, x2, x3;
	output f1, f2;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314, d315, d316, d317, d318, d319, d320, d321, d322, d323, d324, d325, d326, d327, d328, d329, d330, d331, d332, d333, d334, d335, d336, d337, d338, d339, d340, d341, d342, d343, d344, d345, d346, d347, d348, d349, d350, d351, d352, d353, d354, d355, d356, d357, d358, d359, d360, d361, d362, d363, d364, d365, d366, d367, d368, d369, d370, d371, d372, d373;

	not (d1, x1);
	or (d2, x0, x2);
	nand (d3, x1, x2);
	buf (d4, x2);
	or (d5, x0, x3);
	xor (d6, x0, x3);
	xnor (d7, x1, x2);
	xnor (d8, x2, x3);
	xnor (d9, x2);
	and (d10, x1, x3);
	and (d11, x2, x3);
	nor (d12, x2, x3);
	or (d13, x0, x2);
	not (d14, x2);
	buf (d15, x3);
	xor (d16, x0, x1);
	or (d17, x1);
	xnor (d18, x3);
	nand (d19, x1, x2);
	and (d20, x0, x2);
	nor (d21, x2);
	xor (d22, x2, x3);
	xor (d23, x3);
	nand (d24, x1);
	not (d25, x0);
	nor (d26, x2, x3);
	buf (d27, x1);
	or (d28, x3);
	or (d29, x2, x3);
	xnor (d30, x0, x3);
	xnor (d31, x0, x1);
	or (d32, x1, x2);
	nand (d33, x0, x3);
	nand (d34, x0);
	nand (d35, x0, x3);
	nor (d36, x1, x3);
	or (d37, x1, x3);
	buf (d38, x0);
	xor (d39, x0, x1);
	and (d40, x0, x3);
	nand (d41, x0, x1);
	and (d42, x2, x3);
	and (d43, x0, x2);
	or (d44, x0);
	and (d45, x3);
	xor (d46, x1, x2);
	and (d47, x1, x3);
	xnor (d48, x2, x3);
	and (d49, x2);
	or (d50, x2);
	xor (d51, x1, x2);
	xor (d52, x2);
	nand (d53, x2);
	nor (d54, x0, x3);
	and (d55, d18, d24);
	nand (d56, d15, d28);
	or (d57, d10, d15);
	nand (d58, d10, d37);
	nor (d59, d43, d48);
	nor (d60, d1, d34);
	or (d61, d33, d38);
	nor (d62, d15, d38);
	and (d63, d45, d52);
	buf (d64, d40);
	xnor (d65, d19, d46);
	xor (d66, d18, d27);
	nand (d67, d7, d26);
	not (d68, d50);
	nor (d69, d12, d28);
	and (d70, d35, d50);
	nor (d71, d11, d31);
	and (d72, d10, d18);
	or (d73, d26, d49);
	xor (d74, d9, d16);
	xor (d75, d10, d44);
	not (d76, d9);
	not (d77, d11);
	nand (d78, d37, d53);
	buf (d79, d1);
	or (d80, d15, d28);
	and (d81, d12, d28);
	or (d82, d13, d19);
	xor (d83, d20, d43);
	xnor (d84, d2, d18);
	buf (d85, d28);
	xnor (d86, d3, d34);
	or (d87, d21, d28);
	and (d88, d21, d45);
	nand (d89, d30, d41);
	xnor (d90, d36, d51);
	nand (d91, d39, d43);
	nand (d92, d9, d53);
	or (d93, d41, d49);
	not (d94, d10);
	not (d95, d5);
	nor (d96, d19, d28);
	xor (d97, d6, d25);
	xnor (d98, d27, d40);
	not (d99, d54);
	nand (d100, d28, d50);
	nor (d101, d10, d53);
	nand (d102, d1, d36);
	xor (d103, d2, d29);
	buf (d104, d46);
	xnor (d105, d8, d24);
	xor (d106, d26, d51);
	nand (d107, d19, d42);
	and (d108, d23, d46);
	nand (d109, d25, d37);
	or (d110, d20, d34);
	not (d111, d29);
	nor (d112, d37, d44);
	xnor (d113, d1, d23);
	or (d114, d12, d18);
	and (d115, d38, d51);
	and (d116, d9, d38);
	buf (d117, d17);
	xnor (d118, d40);
	or (d119, d7, d49);
	xnor (d120, d6, d13);
	or (d121, d27, d33);
	buf (d122, d16);
	nand (d123, d8, d39);
	xor (d124, d32, d35);
	nor (d125, d5, d31);
	buf (d126, d13);
	nor (d127, d30, d34);
	xor (d128, d23, d52);
	or (d129, d28, d35);
	and (d130, d26, d51);
	and (d131, d28, d37);
	and (d132, d93, d116);
	buf (d133, d62);
	not (d134, d63);
	nand (d135, d93);
	buf (d136, d42);
	xnor (d137, d69, d115);
	buf (d138, d122);
	nand (d139, d57, d95);
	not (d140, d82);
	nor (d141, d106, d124);
	buf (d142, d33);
	nand (d143, d92, d113);
	buf (d144, d69);
	nor (d145, d103, d125);
	not (d146, d74);
	nor (d147, d79, d92);
	or (d148, d59, d85);
	nand (d149, d93, d98);
	xor (d150, d91, d125);
	or (d151, d78, d108);
	or (d152, d64, d101);
	and (d153, d95, d115);
	nor (d154, d66, d108);
	xnor (d155, d97, d100);
	buf (d156, d131);
	or (d157, d87, d115);
	nand (d158, d80, d108);
	or (d159, d55, d69);
	xor (d160, d69, d123);
	buf (d161, d124);
	or (d162, d59, d113);
	xnor (d163, d62, d91);
	xnor (d164, d74, d119);
	or (d165, d100, d122);
	buf (d166, d54);
	nor (d167, d86, d128);
	buf (d168, d23);
	buf (d169, d45);
	xor (d170, d81, d94);
	or (d171, d79, d87);
	xnor (d172, d106, d114);
	not (d173, d99);
	buf (d174, d97);
	nor (d175, d69, d117);
	or (d176, d97, d123);
	xnor (d177, d145, d158);
	nand (d178, d148, d155);
	not (d179, d117);
	or (d180, d152, d161);
	not (d181, d2);
	and (d182, d151, d163);
	not (d183, d105);
	nor (d184, d136, d164);
	xnor (d185, d141, d152);
	nor (d186, d151, d154);
	buf (d187, d140);
	buf (d188, d107);
	not (d189, d96);
	not (d190, d55);
	or (d191, d158, d174);
	xnor (d192, d146);
	nand (d193, d133, d174);
	nor (d194, d167, d171);
	xnor (d195, d168, d171);
	nand (d196, d145, d155);
	xor (d197, d158, d174);
	nor (d198, d172, d176);
	not (d199, d176);
	xor (d200, d143, d144);
	nand (d201, d154, d168);
	xor (d202, d174, d175);
	xnor (d203, d145, d176);
	or (d204, d142, d152);
	not (d205, d119);
	nand (d206, d193, d204);
	xor (d207, d177, d203);
	or (d208, d179, d183);
	or (d209, d195, d197);
	xnor (d210, d180, d183);
	nand (d211, d187, d197);
	buf (d212, d9);
	not (d213, d16);
	and (d214, d187, d194);
	and (d215, d184, d197);
	nand (d216, d181, d192);
	and (d217, d183, d184);
	nor (d218, d184, d202);
	nand (d219, d185, d202);
	nand (d220, d185, d199);
	xor (d221, d190, d191);
	buf (d222, d10);
	buf (d223, d29);
	nand (d224, d177, d193);
	nand (d225, d192, d200);
	buf (d226, d95);
	buf (d227, d92);
	nor (d228, d186);
	xor (d229, d179, d180);
	not (d230, d102);
	xnor (d231, d178, d197);
	not (d232, d17);
	and (d233, d182, d190);
	not (d234, d172);
	xnor (d235, d184, d198);
	buf (d236, d152);
	or (d237, d177, d182);
	nand (d238, d177, d198);
	buf (d239, d25);
	or (d240, d179, d196);
	not (d241, d62);
	xnor (d242, d197, d201);
	and (d243, d181, d203);
	nand (d244, d188, d199);
	nor (d245, d186, d203);
	xnor (d246, d178, d183);
	xor (d247, d177, d199);
	not (d248, d72);
	xor (d249, d180, d201);
	or (d250, d184, d200);
	xor (d251, d187, d199);
	buf (d252, d15);
	or (d253, d184, d199);
	nand (d254, d184, d188);
	nor (d255, d190, d191);
	and (d256, d184, d199);
	nand (d257, d178, d183);
	buf (d258, d155);
	and (d259, d179, d203);
	or (d260, d180, d183);
	and (d261, d181, d183);
	xnor (d262, d177, d204);
	xnor (d263, d185, d187);
	nand (d264, d192, d203);
	not (d265, d203);
	buf (d266, d147);
	xnor (d267, d191, d198);
	buf (d268, d56);
	xnor (d269, d183, d186);
	xnor (d270, d193, d204);
	xor (d271, d181, d192);
	xor (d272, d184, d201);
	or (d273, d189, d204);
	not (d274, d23);
	xor (d275, d183, d203);
	xor (d276, d196, d200);
	or (d277, d188, d200);
	nor (d278, d197, d200);
	xor (d279, d181, d187);
	nor (d280, d190, d201);
	and (d281, d177, d184);
	or (d282, d182, d198);
	nand (d283, d207, d220);
	or (d284, d221, d234);
	xor (d285, d254, d271);
	and (d286, d218, d269);
	or (d287, d209, d223);
	xnor (d288, d233, d245);
	nand (d289, d212, d270);
	nor (d290, d205, d276);
	and (d291, d269, d272);
	buf (d292, d230);
	xnor (d293, d206, d265);
	and (d294, d222, d224);
	nor (d295, d240, d260);
	or (d296, d212, d257);
	and (d297, d214, d247);
	nand (d298, d254, d267);
	and (d299, d208, d269);
	and (d300, d229, d258);
	xnor (d301, d245, d270);
	or (d302, d215, d258);
	and (d303, d216, d254);
	xnor (d304, d268, d272);
	buf (d305, d6);
	xnor (d306, d235, d278);
	nand (d307, d271, d273);
	and (d308, d208, d213);
	xnor (d309, d236, d257);
	and (d310, d251, d262);
	nor (d311, d262, d282);
	and (d312, d215, d278);
	xnor (d313, d241, d254);
	or (d314, d224, d242);
	or (d315, d233, d243);
	xor (d316, d253, d272);
	buf (d317, d20);
	nor (d318, d243, d246);
	not (d319, d263);
	buf (d320, d199);
	nor (d321, d233, d235);
	buf (d322, d43);
	not (d323, d95);
	nand (d324, d262, d279);
	nor (d325, d249, d277);
	xnor (d326, d218, d268);
	nand (d327, d227, d282);
	xnor (d328, d248, d256);
	buf (d329, d143);
	xor (d330, d223, d254);
	xnor (d331, d227, d236);
	and (d332, d261, d267);
	xor (d333, d221, d238);
	xor (d334, d208, d249);
	not (d335, d33);
	or (d336, d232, d259);
	or (d337, d257, d267);
	nor (d338, d239, d271);
	xor (d339, d217, d251);
	buf (d340, d178);
	nand (d341, d208, d252);
	nand (d342, d226, d248);
	or (d343, d222, d255);
	nand (d344, d206, d280);
	buf (d345, d270);
	or (d346, d239, d261);
	xor (d347, d236, d250);
	buf (d348, d70);
	xor (d349, d264, d269);
	nand (d350, d228, d280);
	or (d351, d224, d280);
	or (d352, d255, d276);
	nor (d353, d223, d260);
	xnor (d354, d234, d254);
	nor (d355, d255, d280);
	buf (d356, d109);
	xnor (d357, d213, d259);
	not (d358, d19);
	or (d359, d218, d229);
	nand (d360, d232, d247);
	or (d361, d212, d258);
	xnor (d362, d246, d273);
	buf (d363, d269);
	xor (d364, d235, d236);
	or (d365, d256, d282);
	or (d366, d228, d273);
	or (d367, d243, d268);
	nand (d368, d245, d248);
	nor (d369, d283, d285);
	not (d370, d297);
	and (d371, d309, d343);
	nor (d372, d284, d347);
	or (d373, d305, d341);
	assign f1 = d371;
	assign f2 = d372;
endmodule
