module CCGRCG126( x0, x1, x2, x3, x4, f1, f2, f3, f4, f5, f6, f7, f8 );

	input x0, x1, x2, x3, x4;
	output f1, f2, f3, f4, f5, f6, f7, f8;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248;

	not (d1, x0);
	xor (d2, x2, x3);
	or (d3, x0);
	buf (d4, x0);
	xor (d5, x1, x3);
	or (d6, x2, x4);
	xor (d7, x0, x3);
	xnor (d8, x3, x4);
	buf (d9, x2);
	nor (d10, x1, x3);
	and (d11, x1, x3);
	xor (d12, x0, x1);
	nand (d13, x0, x2);
	nor (d14, x2);
	and (d15, x2);
	nand (d16, x1, x2);
	nand (d17, x2, x4);
	or (d18, x1, x3);
	nor (d19, x0, x2);
	nand (d20, x0, x4);
	or (d21, x0, x1);
	nor (d22, x1, x4);
	xor (d23, x0);
	and (d24, x4);
	or (d25, x0, x3);
	or (d26, x2);
	xnor (d27, x1, x3);
	and (d28, x1, x4);
	nor (d29, x3, x4);
	xnor (d30, x1, x3);
	not (d31, x3);
	buf (d32, x1);
	buf (d33, x3);
	not (d34, x4);
	xnor (d35, x0, x1);
	nor (d36, x4);
	and (d37, x1, x4);
	xor (d38, x1, x4);
	or (d39, x0, x4);
	or (d40, x0, x4);
	or (d41, d7, d37);
	not (d42, d4);
	xnor (d43, d15, d40);
	xor (d44, d10, d25);
	nand (d45, d13, d24);
	and (d46, d24, d36);
	not (d47, d14);
	nor (d48, d19, d27);
	not (d49, d33);
	not (d50, d31);
	xnor (d51, d27, d35);
	buf (d52, d31);
	not (d53, d32);
	nor (d54, d14, d27);
	or (d55, d7, d32);
	buf (d56, d30);
	nand (d57, d8);
	not (d58, d21);
	xnor (d59, d16, d19);
	or (d60, d6, d12);
	or (d61, d6, d30);
	xnor (d62, d13, d34);
	not (d63, d22);
	nor (d64, d16, d36);
	xor (d65, d13, d24);
	or (d66, d22, d34);
	or (d67, d12, d13);
	and (d68, d60, d61);
	nor (d69, d62, d67);
	nor (d70, d44, d48);
	xor (d71, d51, d58);
	buf (d72, d52);
	buf (d73, d38);
	not (d74, d52);
	nand (d75, d53, d66);
	or (d76, d44, d55);
	not (d77, d50);
	xnor (d78, d59, d60);
	or (d79, d50, d65);
	xnor (d80, d50, d65);
	xor (d81, d50, d51);
	buf (d82, d17);
	nand (d83, d59, d66);
	xor (d84, d64, d66);
	xor (d85, d52, d53);
	and (d86, d43, d50);
	nand (d87, d53, d56);
	buf (d88, d2);
	not (d89, d53);
	xnor (d90, d53, d65);
	and (d91, d48, d65);
	nand (d92, d54, d64);
	and (d93, d50, d66);
	not (d94, d6);
	nand (d95, d54, d65);
	or (d96, d41);
	or (d97, d48, d58);
	and (d98, d46, d64);
	not (d99, d25);
	nand (d100, d41, d60);
	xor (d101, d46, d59);
	xnor (d102, d44, d62);
	nand (d103, d41, d51);
	xor (d104, d52, d57);
	buf (d105, d45);
	nand (d106, d43, d61);
	buf (d107, d8);
	or (d108, d42, d66);
	not (d109, d26);
	and (d110, d60, d65);
	buf (d111, d35);
	or (d112, d52, d67);
	buf (d113, d48);
	nand (d114, d58, d59);
	and (d115, d43, d64);
	and (d116, d44, d51);
	or (d117, d78, d86);
	and (d118, d90, d112);
	xnor (d119, d84, d85);
	xnor (d120, d95, d99);
	nor (d121, d85, d99);
	or (d122, d97, d101);
	xnor (d123, d87, d92);
	xor (d124, d94, d114);
	nand (d125, d70, d106);
	or (d126, d108, d116);
	and (d127, d77, d115);
	buf (d128, d107);
	xnor (d129, d98, d102);
	xnor (d130, d80, d99);
	nand (d131, d69, d94);
	and (d132, d89, d108);
	buf (d133, d37);
	buf (d134, d69);
	nand (d135, d84, d102);
	xnor (d136, d76, d112);
	buf (d137, d54);
	not (d138, d10);
	nor (d139, d68, d81);
	xnor (d140, d72, d78);
	nand (d141, d79, d89);
	or (d142, d76, d101);
	nor (d143, d98, d102);
	or (d144, d69, d100);
	or (d145, d99, d109);
	not (d146, d74);
	and (d147, d85, d98);
	nand (d148, d80, d109);
	nand (d149, d74, d90);
	buf (d150, d68);
	nand (d151, d78, d98);
	xnor (d152, d84, d107);
	buf (d153, d11);
	or (d154, d88, d113);
	xnor (d155, d96, d106);
	nand (d156, d82, d102);
	nor (d157, d68, d80);
	not (d158, d79);
	or (d159, d88, d115);
	or (d160, d109, d111);
	or (d161, d68, d69);
	xor (d162, d74, d76);
	or (d163, d76, d103);
	nand (d164, d78, d106);
	xor (d165, d78, d83);
	xnor (d166, d68, d93);
	xor (d167, d78, d102);
	xnor (d168, d90, d93);
	xor (d169, d81, d109);
	or (d170, d70, d111);
	nor (d171, d77, d96);
	not (d172, d98);
	xor (d173, d70, d93);
	not (d174, d19);
	nor (d175, d88, d104);
	not (d176, d92);
	nand (d177, d75, d92);
	xor (d178, d85, d99);
	not (d179, d8);
	or (d180, d86, d93);
	nor (d181, d69, d97);
	buf (d182, d46);
	nand (d183, d101, d112);
	or (d184, d74, d103);
	xor (d185, d98, d101);
	nand (d186, d69, d83);
	xnor (d187, d77, d109);
	not (d188, d68);
	buf (d189, d110);
	xnor (d190, d94, d104);
	and (d191, d79, d89);
	nor (d192, d80, d109);
	xor (d193, d150, d155);
	xor (d194, d132, d143);
	and (d195, d152, d186);
	or (d196, d134, d145);
	or (d197, d171, d182);
	xnor (d198, d171, d191);
	or (d199, d162, d178);
	nand (d200, d134, d164);
	nor (d201, d157, d160);
	xnor (d202, d122, d162);
	or (d203, d174, d190);
	nor (d204, d154, d164);
	or (d205, d135, d164);
	nor (d206, d177, d179);
	buf (d207, d138);
	and (d208, d135, d183);
	xnor (d209, d147, d180);
	and (d210, d148, d186);
	buf (d211, d58);
	xnor (d212, d156, d160);
	nand (d213, d120, d168);
	and (d214, d155, d177);
	buf (d215, d167);
	xnor (d216, d119, d161);
	xnor (d217, d119, d124);
	buf (d218, d114);
	and (d219, d124, d144);
	not (d220, d143);
	xnor (d221, d130, d141);
	nor (d222, d123, d150);
	nand (d223, d157, d175);
	xnor (d224, d118, d150);
	nor (d225, d150, d171);
	and (d226, d161, d177);
	nor (d227, d123, d148);
	and (d228, d122, d134);
	xor (d229, d141, d191);
	or (d230, d144, d152);
	and (d231, d183, d191);
	nand (d232, d128, d164);
	not (d233, d162);
	nand (d234, d137, d186);
	and (d235, d142, d161);
	and (d236, d164, d183);
	or (d237, d118, d181);
	not (d238, d190);
	xor (d239, d154, d183);
	xnor (d240, d151, d154);
	not (d241, d146);
	nand (d242, d174, d187);
	or (d243, d139, d158);
	xnor (d244, d128, d151);
	or (d245, d133, d168);
	xnor (d246, d168, d171);
	nand (d247, d134, d165);
	and (d248, d131, d141);
	assign f1 = d195;
	assign f2 = d224;
	assign f3 = d231;
	assign f4 = d212;
	assign f5 = d210;
	assign f6 = d230;
	assign f7 = d220;
	assign f8 = d244;
endmodule
