module CCGRCG200( x0, x1, x2, x3, x4, x5, x6, f1, f2, f3, f4, f5, f6, f7 );

	input x0, x1, x2, x3, x4, x5, x6;
	output f1, f2, f3, f4, f5, f6, f7;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314, d315, d316, d317, d318, d319, d320, d321, d322;

	nor (d1, x0, x4);
	or (d2, x3, x6);
	xor (d3, x0, x2);
	buf (d4, x6);
	nand (d5, x1, x3);
	not (d6, x1);
	xnor (d7, x3, x4);
	xor (d8, x2, x6);
	nand (d9, x0, x5);
	buf (d10, x3);
	nor (d11, x0, x4);
	nor (d12, x1, x5);
	nor (d13, x3, x6);
	xor (d14, x2, x5);
	nand (d15, x2, x6);
	and (d16, x1, x2);
	not (d17, x2);
	not (d18, x4);
	buf (d19, x5);
	buf (d20, x2);
	buf (d21, x4);
	nand (d22, x0, x3);
	or (d23, x3);
	and (d24, x4, x6);
	nand (d25, x0, x4);
	nor (d26, x0);
	not (d27, x3);
	xor (d28, x1, x3);
	nor (d29, d10, d28);
	nand (d30, d3);
	nand (d31, d2, d11);
	buf (d32, d28);
	nor (d33, d2, d4);
	xnor (d34, d16, d19);
	or (d35, d7, d17);
	xnor (d36, d8, d16);
	nor (d37, d9, d16);
	xor (d38, d1, d21);
	nor (d39, d13, d23);
	xor (d40, d23, d25);
	xnor (d41, d25, d28);
	xnor (d42, d9, d14);
	or (d43, d3, d22);
	xor (d44, d11, d15);
	nor (d45, d5, d23);
	not (d46, d25);
	not (d47, d28);
	nand (d48, d14);
	not (d49, d2);
	xor (d50, d3, d18);
	nand (d51, d23, d27);
	xnor (d52, d2, d18);
	buf (d53, d18);
	nand (d54, d3, d20);
	nand (d55, d1, d25);
	and (d56, d2, d18);
	not (d57, d9);
	and (d58, d1, d6);
	nor (d59, d1, d4);
	nor (d60, d9, d14);
	not (d61, d11);
	or (d62, d14, d16);
	nand (d63, d17, d24);
	xor (d64, d2, d27);
	nor (d65, d12);
	xor (d66, d7, d14);
	not (d67, d26);
	and (d68, d4, d8);
	or (d69, d9, d16);
	xnor (d70, d2, d11);
	nor (d71, d14, d19);
	nor (d72, d2, d16);
	xor (d73, d12, d23);
	or (d74, d24, d27);
	xnor (d75, d18, d27);
	not (d76, d22);
	not (d77, d7);
	and (d78, d15, d21);
	xor (d79, d7, d28);
	and (d80, d8, d25);
	and (d81, d7, d13);
	or (d82, d7, d15);
	xnor (d83, d1, d18);
	nor (d84, d12, d27);
	or (d85, d2, d4);
	nor (d86, d17, d18);
	and (d87, d6, d27);
	and (d88, d24, d26);
	xnor (d89, d9, d18);
	nand (d90, d10, d19);
	and (d91, d20, d24);
	and (d92, d44, d46);
	and (d93, d61, d62);
	buf (d94, d47);
	xnor (d95, d39, d58);
	xnor (d96, d34, d64);
	nand (d97, d32, d90);
	and (d98, d66, d68);
	or (d99, d76, d80);
	nand (d100, d49, d76);
	not (d101, d35);
	buf (d102, d41);
	nor (d103, d63, d64);
	and (d104, d34, d69);
	buf (d105, d17);
	buf (d106, d27);
	xnor (d107, d35, d53);
	buf (d108, d21);
	nor (d109, d53, d68);
	nor (d110, d42, d64);
	nand (d111, d42, d45);
	and (d112, d29, d34);
	or (d113, d32, d80);
	buf (d114, d19);
	nor (d115, d31, d64);
	not (d116, d62);
	nand (d117, d31, d42);
	not (d118, d57);
	or (d119, d34, d91);
	and (d120, d50, d84);
	xor (d121, d38, d76);
	xor (d122, d33, d90);
	xor (d123, d37, d79);
	or (d124, d65, d83);
	or (d125, d39, d82);
	nand (d126, d38, d78);
	xnor (d127, d33, d45);
	or (d128, d69, d87);
	nor (d129, d63, d85);
	nor (d130, d55, d82);
	buf (d131, d72);
	nand (d132, d50, d51);
	nand (d133, d35, d91);
	nand (d134, d45, d59);
	and (d135, d30, d49);
	nand (d136, d30, d85);
	xnor (d137, d34, d35);
	nand (d138, d30, d53);
	nor (d139, d50, d64);
	xor (d140, d64, d82);
	buf (d141, d48);
	nor (d142, d60, d90);
	nor (d143, d38, d67);
	buf (d144, d26);
	xor (d145, d38, d75);
	xnor (d146, d43, d50);
	buf (d147, d59);
	and (d148, d36, d73);
	nor (d149, d49, d87);
	xor (d150, d41, d59);
	or (d151, d39, d74);
	and (d152, d45, d72);
	nor (d153, d31, d38);
	xnor (d154, d58, d68);
	buf (d155, d69);
	nor (d156, d33, d58);
	not (d157, d68);
	nand (d158, d42, d80);
	nor (d159, d59, d79);
	xnor (d160, d80, d89);
	buf (d161, d77);
	buf (d162, d10);
	nor (d163, d49, d65);
	xor (d164, d56, d60);
	xnor (d165, d33, d74);
	nand (d166, d29, d67);
	xor (d167, d76, d78);
	buf (d168, d35);
	xnor (d169, d45, d91);
	or (d170, d35, d69);
	buf (d171, d70);
	xnor (d172, d58, d73);
	nor (d173, d33, d53);
	not (d174, d20);
	and (d175, d66, d83);
	xnor (d176, d39, d44);
	buf (d177, d86);
	xor (d178, d48, d50);
	not (d179, d84);
	and (d180, d60, d68);
	buf (d181, d81);
	nand (d182, d71, d75);
	xnor (d183, d38, d57);
	nand (d184, d51, d76);
	nand (d185, d104, d174);
	or (d186, d126, d141);
	nand (d187, d127, d177);
	buf (d188, d4);
	nand (d189, d123, d152);
	xnor (d190, d101, d107);
	and (d191, d110, d144);
	xor (d192, d94, d135);
	nand (d193, d141, d182);
	not (d194, d138);
	nor (d195, d102, d158);
	or (d196, d96, d153);
	xnor (d197, d137, d173);
	xnor (d198, d108, d118);
	buf (d199, d42);
	nand (d200, d138, d159);
	and (d201, d142, d155);
	not (d202, d135);
	not (d203, d19);
	and (d204, d111, d173);
	xor (d205, d144, d182);
	nand (d206, d157, d158);
	buf (d207, d156);
	and (d208, d110, d173);
	xor (d209, d118, d173);
	nor (d210, d104, d135);
	nor (d211, d113, d126);
	nand (d212, d126, d142);
	nor (d213, d93, d158);
	nand (d214, d136, d178);
	or (d215, d131, d179);
	or (d216, d130, d140);
	xor (d217, d148, d154);
	xor (d218, d112, d157);
	xnor (d219, d96, d119);
	buf (d220, d68);
	xnor (d221, d121, d159);
	xor (d222, d124, d139);
	xnor (d223, d96, d175);
	xor (d224, d161, d162);
	or (d225, d146, d178);
	not (d226, d59);
	buf (d227, d90);
	xor (d228, d152, d171);
	xnor (d229, d117, d119);
	xnor (d230, d203, d228);
	or (d231, d203, d217);
	nand (d232, d224, d225);
	or (d233, d200, d210);
	and (d234, d192, d218);
	nor (d235, d201, d206);
	buf (d236, d71);
	and (d237, d194, d201);
	nand (d238, d204, d219);
	and (d239, d187, d191);
	xnor (d240, d220, d229);
	xnor (d241, d198, d225);
	or (d242, d191, d226);
	not (d243, d156);
	nand (d244, d203, d216);
	xor (d245, d185, d199);
	not (d246, d14);
	nor (d247, d216, d221);
	nor (d248, d209, d222);
	or (d249, d186, d213);
	not (d250, d198);
	nand (d251, d209, d214);
	xnor (d252, d185, d219);
	or (d253, d187);
	nand (d254, d205, d208);
	nand (d255, d212, d219);
	buf (d256, d192);
	nand (d257, d211, d212);
	nand (d258, d222, d225);
	buf (d259, d167);
	or (d260, d199, d229);
	xor (d261, d200, d201);
	not (d262, d115);
	xor (d263, d208, d229);
	nor (d264, d196, d225);
	buf (d265, d97);
	and (d266, d211, d216);
	nand (d267, d188, d228);
	buf (d268, d111);
	nand (d269, d191, d195);
	xor (d270, d188, d227);
	xor (d271, d190, d229);
	buf (d272, d104);
	or (d273, d193, d207);
	nand (d274, d185, d197);
	nor (d275, d201, d210);
	xor (d276, d208, d221);
	or (d277, d189, d224);
	nor (d278, d186, d218);
	and (d279, d200, d215);
	xor (d280, d202, d228);
	nor (d281, d195, d205);
	buf (d282, d55);
	buf (d283, d136);
	nand (d284, d191, d193);
	xor (d285, d189, d209);
	nor (d286, d214, d227);
	xnor (d287, d194, d225);
	xor (d288, d194, d220);
	xnor (d289, d188, d190);
	or (d290, d210, d227);
	not (d291, d216);
	and (d292, d194, d219);
	nor (d293, d200, d218);
	nor (d294, d187, d205);
	buf (d295, d14);
	nor (d296, d199, d221);
	nand (d297, d191, d204);
	xor (d298, d185, d203);
	nand (d299, d210, d225);
	xor (d300, d201, d229);
	xor (d301, d199, d204);
	and (d302, d207, d219);
	buf (d303, d181);
	or (d304, d194, d195);
	not (d305, x0);
	nand (d306, d203, d216);
	nand (d307, d205, d217);
	xnor (d308, d199, d210);
	buf (d309, d13);
	xnor (d310, d191, d224);
	xnor (d311, d188, d192);
	nand (d312, d193, d206);
	not (d313, d158);
	and (d314, d190, d218);
	xor (d315, d204, d226);
	and (d316, d203, d227);
	nand (d317, d188, d214);
	and (d318, d201, d207);
	or (d319, d193, d215);
	nor (d320, d192, d206);
	nor (d321, d199, d223);
	xnor (d322, d203, d219);
	assign f1 = d268;
	assign f2 = d310;
	assign f3 = d297;
	assign f4 = d241;
	assign f5 = d277;
	assign f6 = d319;
	assign f7 = d285;
endmodule
