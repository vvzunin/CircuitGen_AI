module CCGRCG92( x0, x1, x2, x3, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10 );

	input x0, x1, x2, x3;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133;

	nor (d1, x0, x3);
	or (d2, x0, x3);
	and (d3, x0, x2);
	and (d4, x3);
	buf (d5, x1);
	nand (d6, x0, x2);
	nand (d7, x0, x1);
	nor (d8, x1);
	nor (d9, x0, x1);
	nand (d10, x0, x2);
	xnor (d11, x0, x1);
	not (d12, x1);
	nor (d13, x0);
	nor (d14, x2, x3);
	xnor (d15, x2, x3);
	and (d16, x0, x1);
	or (d17, x0);
	nand (d18, x3);
	xor (d19, x0);
	buf (d20, x3);
	nand (d21, x1);
	and (d22, x1, x2);
	nand (d23, x1, x3);
	not (d24, x3);
	xnor (d25, x0);
	and (d26, x1, x2);
	or (d27, x1, x2);
	xor (d28, x1, x2);
	and (d29, x2);
	and (d30, x0, x3);
	not (d31, x0);
	xnor (d32, x1, x2);
	nor (d33, x0, x3);
	nand (d34, x0, x3);
	and (d35, x2, x3);
	or (d36, x1, x3);
	or (d37, x0, x3);
	and (d38, x0, x1);
	not (d39, x2);
	nor (d40, x2, x3);
	xnor (d41, x0, x2);
	xor (d42, x0, x3);
	or (d43, x3);
	xor (d44, x0, x1);
	buf (d45, x2);
	xor (d46, x0, x1);
	xor (d47, x0, x2);
	xor (d48, x1, x3);
	nand (d49, x0, x3);
	xor (d50, x2, x3);
	and (d51, x2, x3);
	or (d52, x2, x3);
	or (d53, x2);
	and (d54, x1, x3);
	nand (d55, x1, x2);
	nand (d56, x0, x1);
	xor (d57, x0, x2);
	xnor (d58, x1);
	nor (d59, x1, x3);
	buf (d60, d6);
	nand (d61, d23, d49);
	nand (d62, d9, d34);
	not (d63, d50);
	buf (d64, d37);
	not (d65, d45);
	nor (d66, d44, d56);
	nand (d67, d37, d53);
	nor (d68, d16, d45);
	or (d69, d2, d57);
	not (d70, d5);
	and (d71, d45, d55);
	nand (d72, d2, d54);
	buf (d73, d21);
	xor (d74, d18, d23);
	nor (d75, d13, d47);
	xnor (d76, d8, d16);
	nand (d77, d19, d57);
	or (d78, d16, d59);
	nand (d79, d11, d54);
	buf (d80, d23);
	nand (d81, d32, d44);
	nand (d82, d9, d48);
	nor (d83, d7, d32);
	xnor (d84, d35, d43);
	xor (d85, d44, d57);
	nand (d86, d13, d37);
	xnor (d87, d1, d11);
	or (d88, d29, d53);
	or (d89, d6, d20);
	or (d90, d10, d34);
	nand (d91, d32, d40);
	xor (d92, d36, d41);
	nor (d93, d58, d59);
	xor (d94, d18, d34);
	xor (d95, d9, d58);
	and (d96, d13, d55);
	nand (d97, d51, d58);
	buf (d98, d45);
	nand (d99, d33, d49);
	or (d100, d2, d59);
	not (d101, d13);
	or (d102, d30, d48);
	nor (d103, d22, d27);
	nand (d104, d2, d59);
	xnor (d105, d1, d52);
	xor (d106, d28, d58);
	xnor (d107, d5, d40);
	buf (d108, d30);
	nand (d109, d2, d13);
	or (d110, d12, d44);
	nor (d111, d27, d36);
	nand (d112, d10, d36);
	and (d113, d6, d13);
	or (d114, d21, d39);
	and (d115, d19, d39);
	nand (d116, d11, d22);
	buf (d117, d50);
	xnor (d118, d48, d58);
	nor (d119, d29, d54);
	xor (d120, d4, d54);
	buf (d121, d43);
	and (d122, d5, d45);
	nand (d123, d14, d46);
	and (d124, d18, d33);
	xor (d125, d43, d50);
	xnor (d126, d8, d17);
	not (d127, d24);
	xor (d128, d3, d51);
	or (d129, d14, d57);
	xnor (d130, d32, d47);
	not (d131, d19);
	not (d132, d52);
	xor (d133, d25, d37);
	assign f1 = d66;
	assign f2 = d112;
	assign f3 = d63;
	assign f4 = d129;
	assign f5 = d115;
	assign f6 = d78;
	assign f7 = d122;
	assign f8 = d104;
	assign f9 = d129;
	assign f10 = d84;
endmodule
