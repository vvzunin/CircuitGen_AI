module CCGRCG134( x0, x1, x2, x3, x4, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12 );

	input x0, x1, x2, x3, x4;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261;

	xor (d1, x0, x3);
	and (d2, x2, x3);
	buf (d3, x3);
	and (d4, x0, x1);
	nand (d5, x1, x3);
	and (d6, x1, x4);
	nor (d7, x1);
	not (d8, x2);
	nand (d9, x0, x1);
	buf (d10, x0);
	buf (d11, x2);
	buf (d12, x4);
	or (d13, x1, x3);
	and (d14, x0, x3);
	not (d15, x4);
	nand (d16, x2);
	not (d17, x1);
	nand (d18, x0, x2);
	xnor (d19, x1, x4);
	xor (d20, x4);
	nor (d21, x1, x4);
	or (d22, x4);
	xnor (d23, x2, x3);
	or (d24, x1, x4);
	and (d25, x0, x2);
	buf (d26, x1);
	nand (d27, x1, x4);
	nor (d28, x0, x2);
	xor (d29, x0, x3);
	nand (d30, x0, x2);
	xor (d31, x0, x4);
	or (d32, x2);
	xnor (d33, x0, x3);
	xor (d34, x1, x4);
	not (d35, x3);
	nand (d36, x0, x3);
	nand (d37, x2, x3);
	nand (d38, x0, x4);
	or (d39, x2, x4);
	xnor (d40, x0, x4);
	nor (d41, x2, x3);
	or (d42, x0);
	nand (d43, x0);
	nand (d44, x0, x4);
	nor (d45, x2, x4);
	not (d46, x0);
	xor (d47, x1);
	or (d48, x3, x4);
	nor (d49, d21, d39);
	nor (d50, d32, d48);
	and (d51, d5, d8);
	xor (d52, d5, d15);
	xor (d53, d11, d21);
	nor (d54, d1, d31);
	xnor (d55, d33, d44);
	or (d56, d2);
	xnor (d57, d2, d13);
	buf (d58, d7);
	or (d59, d12, d17);
	and (d60, d42, d45);
	nor (d61, d26, d29);
	buf (d62, d8);
	not (d63, d10);
	and (d64, d10, d12);
	xnor (d65, d13, d26);
	xnor (d66, d14, d29);
	not (d67, d14);
	buf (d68, d23);
	or (d69, d1, d3);
	xor (d70, d1, d20);
	or (d71, d32, d34);
	xor (d72, d37, d41);
	nand (d73, d10, d12);
	and (d74, d6, d19);
	nand (d75, d1, d16);
	nand (d76, d9, d33);
	xnor (d77, d31, d35);
	or (d78, d10, d41);
	and (d79, d12, d22);
	and (d80, d35, d43);
	or (d81, d14, d34);
	xnor (d82, d33);
	or (d83, d13, d42);
	xor (d84, d18, d20);
	and (d85, d6, d23);
	xor (d86, d6, d23);
	and (d87, d3, d27);
	nand (d88, d40, d44);
	and (d89, d37, d41);
	and (d90, d6, d32);
	not (d91, d34);
	and (d92, d33, d44);
	buf (d93, d46);
	or (d94, d27, d43);
	not (d95, d29);
	nor (d96, d16, d28);
	nand (d97, d2, d6);
	or (d98, d30, d46);
	and (d99, d17, d30);
	nor (d100, d3, d4);
	and (d101, d51, d64);
	not (d102, d47);
	nand (d103, d93, d96);
	and (d104, d67, d100);
	xnor (d105, d77, d83);
	nor (d106, d77, d79);
	or (d107, d69, d81);
	and (d108, d59, d85);
	nor (d109, d62, d69);
	nor (d110, d56, d72);
	or (d111, d70, d86);
	or (d112, d61, d63);
	or (d113, d88, d97);
	buf (d114, d6);
	nand (d115, d53, d67);
	nor (d116, d52, d89);
	and (d117, d72, d100);
	and (d118, d62, d93);
	xor (d119, d63, d79);
	and (d120, d58, d82);
	nand (d121, d55, d68);
	not (d122, d80);
	and (d123, d74, d85);
	nor (d124, d80, d97);
	or (d125, d56, d63);
	not (d126, d68);
	not (d127, d25);
	not (d128, d35);
	or (d129, d85, d89);
	buf (d130, d9);
	buf (d131, d88);
	nand (d132, d90, d95);
	xnor (d133, d83, d90);
	buf (d134, d50);
	xor (d135, d51, d84);
	or (d136, d67, d75);
	nand (d137, d74, d99);
	buf (d138, d35);
	xnor (d139, d53, d62);
	xor (d140, d61, d98);
	or (d141, d86, d95);
	nor (d142, d50, d58);
	not (d143, d15);
	xnor (d144, d67, d83);
	or (d145, d74, d77);
	not (d146, d20);
	xor (d147, d76, d93);
	nor (d148, d55, d81);
	not (d149, d79);
	and (d150, d66, d84);
	not (d151, d32);
	xor (d152, d57, d63);
	nor (d153, d53, d97);
	buf (d154, d71);
	not (d155, d82);
	or (d156, d134, d147);
	not (d157, d114);
	and (d158, d125, d140);
	xnor (d159, d124, d149);
	and (d160, d114, d149);
	buf (d161, d15);
	xor (d162, d124, d153);
	buf (d163, d41);
	xnor (d164, d125, d128);
	xor (d165, d130, d147);
	nand (d166, d113, d151);
	xor (d167, d133, d153);
	not (d168, d75);
	nand (d169, d122, d152);
	nor (d170, d127, d138);
	xnor (d171, d105, d138);
	or (d172, d131, d154);
	not (d173, d115);
	nand (d174, d132, d137);
	xnor (d175, d116, d139);
	xor (d176, d131, d145);
	xnor (d177, d140, d153);
	not (d178, d81);
	xnor (d179, d102, d108);
	xnor (d180, d106, d114);
	nor (d181, d117, d129);
	or (d182, d114, d141);
	and (d183, d107, d115);
	buf (d184, d62);
	nand (d185, d129, d152);
	xor (d186, d107, d122);
	nand (d187, d126, d154);
	and (d188, d104, d125);
	and (d189, d120, d141);
	not (d190, d18);
	and (d191, d137, d151);
	buf (d192, d95);
	buf (d193, d100);
	nor (d194, d134, d137);
	nor (d195, d130, d152);
	nor (d196, d163, d192);
	xor (d197, d169, d195);
	and (d198, d186, d187);
	buf (d199, d86);
	xnor (d200, d163, d192);
	xnor (d201, d162, d184);
	not (d202, d4);
	xnor (d203, d165, d167);
	and (d204, d200, d202);
	buf (d205, d169);
	buf (d206, d102);
	xor (d207, d197, d198);
	and (d208, d199);
	xor (d209, d199, d202);
	buf (d210, d54);
	nand (d211, d200, d201);
	not (d212, d42);
	and (d213, d197, d199);
	buf (d214, d1);
	nand (d215, d198, d200);
	nor (d216, d196, d201);
	xor (d217, d198, d203);
	xnor (d218, d196, d203);
	xor (d219, d197, d202);
	xnor (d220, d196, d197);
	xnor (d221, d196, d200);
	xnor (d222, d198, d203);
	buf (d223, d158);
	buf (d224, d68);
	xor (d225, d196);
	xnor (d226, d198);
	not (d227, d76);
	or (d228, d197, d201);
	xnor (d229, d197, d203);
	or (d230, d200, d202);
	buf (d231, d164);
	buf (d232, d81);
	and (d233, d196);
	or (d234, d201);
	or (d235, d196, d198);
	xor (d236, d199);
	and (d237, d202);
	nand (d238, d196, d203);
	and (d239, d201);
	and (d240, d202, d203);
	xor (d241, d197, d203);
	or (d242, d197, d198);
	xor (d243, d200, d202);
	and (d244, d198, d203);
	or (d245, d201, d202);
	xnor (d246, d197, d202);
	xor (d247, d196, d200);
	not (d248, d88);
	buf (d249, d179);
	nand (d250, d196);
	nor (d251, d202);
	nor (d252, d197, d202);
	not (d253, d3);
	not (d254, d43);
	not (d255, d12);
	nor (d256, d196, d198);
	nor (d257, d201, d202);
	xnor (d258, d196, d201);
	and (d259, d198, d200);
	xnor (d260, d199, d201);
	and (d261, d198, d202);
	assign f1 = d245;
	assign f2 = d227;
	assign f3 = d252;
	assign f4 = d240;
	assign f5 = d225;
	assign f6 = d227;
	assign f7 = d208;
	assign f8 = d205;
	assign f9 = d223;
	assign f10 = d205;
	assign f11 = d260;
	assign f12 = d211;
endmodule
