module CCGRCG127( x0, x1, x2, x3, x4, f1, f2, f3, f4, f5, f6, f7, f8 );

	input x0, x1, x2, x3, x4;
	output f1, f2, f3, f4, f5, f6, f7, f8;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314, d315, d316, d317, d318, d319, d320, d321, d322, d323, d324, d325, d326, d327, d328, d329, d330, d331, d332, d333, d334, d335, d336, d337, d338, d339, d340, d341, d342, d343, d344, d345, d346, d347, d348, d349, d350, d351, d352, d353, d354, d355, d356, d357, d358, d359, d360, d361, d362, d363, d364, d365, d366, d367, d368, d369, d370, d371, d372, d373, d374, d375, d376, d377, d378, d379, d380, d381, d382, d383, d384, d385, d386, d387, d388, d389, d390, d391, d392, d393, d394, d395, d396, d397, d398, d399, d400, d401, d402, d403, d404, d405, d406, d407, d408, d409, d410, d411, d412, d413, d414, d415, d416, d417, d418, d419, d420, d421, d422, d423;

	buf (d1, x2);
	or (d2, x1, x4);
	not (d3, x3);
	xnor (d4, x2);
	buf (d5, x1);
	nor (d6, x0, x3);
	xor (d7, x0, x1);
	xnor (d8, x0, x1);
	or (d9, x2);
	xor (d10, x2);
	and (d11, x0, x3);
	xnor (d12, x1, x4);
	not (d13, x2);
	not (d14, x0);
	xnor (d15, x2, x4);
	nor (d16, x2, x4);
	xnor (d17, x0, x4);
	nor (d18, x2, x3);
	xor (d19, x0, x4);
	xor (d20, x1, x2);
	buf (d21, x4);
	nand (d22, x0, x4);
	xnor (d23, x0, x2);
	xnor (d24, x4);
	or (d25, x3, x4);
	xor (d26, x0, x4);
	nor (d27, x3);
	not (d28, x1);
	xor (d29, x1, x3);
	or (d30, x1);
	xor (d31, x2, x4);
	nor (d32, x2, x4);
	nand (d33, x0, x1);
	nor (d34, d14, d33);
	or (d35, d16, d27);
	xnor (d36, d15, d30);
	buf (d37, d11);
	nor (d38, d9, d17);
	nand (d39, d1, d32);
	nor (d40, d9, d13);
	not (d41, d11);
	or (d42, d16, d33);
	not (d43, d14);
	xor (d44, d28, d32);
	or (d45, d2, d26);
	and (d46, d4, d30);
	buf (d47, d29);
	xor (d48, d19, d27);
	nand (d49, d5, d17);
	xor (d50, d27, d32);
	not (d51, d1);
	or (d52, d4, d13);
	buf (d53, d22);
	nor (d54, d8, d10);
	nor (d55, d6, d7);
	not (d56, d6);
	nor (d57, d13, d21);
	not (d58, d5);
	xor (d59, d9, d31);
	xnor (d60, d30, d32);
	buf (d61, d14);
	nand (d62, d6, d12);
	buf (d63, d5);
	nand (d64, d10, d13);
	and (d65, d22, d31);
	not (d66, d17);
	buf (d67, d4);
	nand (d68, d5, d9);
	or (d69, d9, d21);
	buf (d70, d23);
	xor (d71, d6, d14);
	buf (d72, d12);
	or (d73, d21, d29);
	xor (d74, d2, d6);
	or (d75, d12, d33);
	xnor (d76, d8, d33);
	xnor (d77, d5);
	buf (d78, d25);
	not (d79, d29);
	not (d80, d23);
	or (d81, d12, d13);
	nor (d82, d1, d8);
	nor (d83, d4, d31);
	nor (d84, d13, d22);
	xor (d85, d8, d17);
	not (d86, d13);
	or (d87, d31);
	nand (d88, d51, d58);
	and (d89, d57, d83);
	xnor (d90, d53, d84);
	xor (d91, d39, d67);
	buf (d92, d36);
	buf (d93, d33);
	or (d94, d52, d71);
	and (d95, d41, d74);
	nor (d96, d48, d54);
	nand (d97, d61, d74);
	and (d98, d59, d64);
	xnor (d99, d39, d87);
	xnor (d100, d52);
	buf (d101, d21);
	buf (d102, d45);
	buf (d103, d48);
	nand (d104, d36, d40);
	xor (d105, d34, d64);
	xor (d106, d66, d86);
	not (d107, d58);
	nor (d108, d34, d37);
	xor (d109, d38, d83);
	or (d110, d68, d70);
	and (d111, d53, d76);
	not (d112, d9);
	xnor (d113, d54, d77);
	not (d114, d40);
	xnor (d115, d39, d43);
	xor (d116, d42, d61);
	or (d117, d111, d113);
	nand (d118, d98, d103);
	not (d119, x4);
	and (d120, d106, d113);
	xnor (d121, d104, d110);
	nand (d122, d99, d113);
	xnor (d123, d105, d111);
	xnor (d124, d102, d104);
	nor (d125, d107, d108);
	or (d126, d114, d116);
	nand (d127, d97, d114);
	and (d128, d91, d97);
	or (d129, d98, d116);
	nor (d130, d95, d96);
	xor (d131, d93, d99);
	nand (d132, d112, d114);
	or (d133, d90, d109);
	not (d134, d75);
	not (d135, d34);
	xnor (d136, d111);
	xor (d137, d91, d113);
	xor (d138, d99, d108);
	and (d139, d97, d112);
	xor (d140, d103, d106);
	xor (d141, d93, d104);
	not (d142, d70);
	and (d143, d90, d114);
	xor (d144, d101, d105);
	and (d145, d103, d108);
	xnor (d146, d106, d109);
	not (d147, d100);
	xnor (d148, d101, d106);
	nor (d149, d98, d112);
	xnor (d150, d95, d116);
	or (d151, d109, d113);
	xnor (d152, d89, d115);
	not (d153, d50);
	buf (d154, d13);
	or (d155, d92, d99);
	not (d156, d84);
	nand (d157, d100, d114);
	or (d158, d100, d101);
	nand (d159, d95, d106);
	buf (d160, d99);
	xor (d161, d103, d111);
	nor (d162, d97, d109);
	or (d163, d103, d110);
	not (d164, d59);
	not (d165, d71);
	xnor (d166, d98, d115);
	not (d167, d10);
	and (d168, d96, d115);
	buf (d169, d19);
	or (d170, d91, d103);
	nor (d171, d93, d97);
	nor (d172, d110, d115);
	and (d173, d91, d107);
	and (d174, d92, d102);
	and (d175, d115);
	nand (d176, d99, d108);
	nor (d177, d96, d115);
	buf (d178, d56);
	buf (d179, d15);
	nand (d180, d103, d110);
	nor (d181, d95, d99);
	not (d182, d56);
	not (d183, d66);
	and (d184, d100, d105);
	nand (d185, d101, d107);
	and (d186, d103, d111);
	or (d187, d112, d116);
	nand (d188, d88, d95);
	xor (d189, d99, d116);
	xor (d190, d92, d97);
	xnor (d191, d89, d90);
	not (d192, d68);
	buf (d193, d103);
	and (d194, d95, d116);
	not (d195, d97);
	nand (d196, d100, d102);
	not (d197, d32);
	and (d198, d109, d110);
	or (d199, d102, d114);
	xor (d200, d91, d97);
	or (d201, d104, d110);
	nand (d202, d90, d100);
	xnor (d203, d102, d107);
	nand (d204, d97, d115);
	nand (d205, d109, d112);
	and (d206, d95, d96);
	xor (d207, d111, d116);
	or (d208, d99, d115);
	xnor (d209, d109, d112);
	not (d210, d35);
	xor (d211, d91, d111);
	xor (d212, d89, d116);
	nand (d213, d142, d176);
	and (d214, d132, d158);
	buf (d215, d106);
	xnor (d216, d127, d163);
	and (d217, d136, d146);
	not (d218, d24);
	not (d219, d102);
	or (d220, d132, d154);
	xnor (d221, d130, d170);
	and (d222, d139, d192);
	and (d223, d186, d206);
	buf (d224, d130);
	and (d225, d157, d162);
	nand (d226, d131, d139);
	nand (d227, d126, d205);
	or (d228, d119, d158);
	buf (d229, d183);
	nand (d230, d164, d168);
	nor (d231, d125, d171);
	and (d232, d169, d192);
	and (d233, d219, d224);
	and (d234, d224, d229);
	nand (d235, d223, d225);
	or (d236, d224, d227);
	or (d237, d218, d219);
	or (d238, d221, d224);
	and (d239, d220, d227);
	and (d240, d218, d224);
	xor (d241, d225, d226);
	buf (d242, d151);
	or (d243, d220, d230);
	xnor (d244, d213, d229);
	not (d245, d162);
	xnor (d246, d215, d226);
	buf (d247, d229);
	xor (d248, d223, d230);
	nor (d249, d218, d219);
	xnor (d250, d228, d232);
	nand (d251, d222, d227);
	not (d252, d152);
	xor (d253, d218, d228);
	nor (d254, d214, d230);
	and (d255, d218, d220);
	nor (d256, d222, d230);
	xnor (d257, d226, d232);
	xor (d258, d223, d230);
	not (d259, d199);
	or (d260, d221, d230);
	not (d261, d103);
	xnor (d262, d218, d227);
	nor (d263, d215, d222);
	not (d264, d36);
	nor (d265, d228, d232);
	and (d266, d216, d223);
	xnor (d267, d216, d217);
	not (d268, d101);
	nand (d269, d219, d220);
	xor (d270, d213, d220);
	and (d271, d222, d231);
	xor (d272, d217, d224);
	nor (d273, d220, d230);
	xnor (d274, d225, d228);
	buf (d275, d105);
	and (d276, d221, d228);
	xnor (d277, d220, d228);
	xor (d278, d218, d226);
	xnor (d279, d215, d228);
	buf (d280, d143);
	buf (d281, d77);
	nand (d282, d225, d228);
	not (d283, d218);
	not (d284, d113);
	and (d285, d219, d230);
	not (d286, d148);
	and (d287, d218, d224);
	nor (d288, d216, d229);
	xnor (d289, d224, d232);
	or (d290, d225, d227);
	xnor (d291, d219, d232);
	xor (d292, d226, d230);
	or (d293, d218);
	and (d294, d219, d229);
	nor (d295, d217, d218);
	not (d296, d2);
	nor (d297, d225, d226);
	or (d298, d213, d216);
	nor (d299, d222);
	buf (d300, d220);
	nor (d301, d216, d226);
	not (d302, d65);
	not (d303, d232);
	xor (d304, d223, d226);
	buf (d305, d224);
	nor (d306, d213, d215);
	buf (d307, d165);
	or (d308, d220, d224);
	nor (d309, d220, d226);
	and (d310, d225, d232);
	and (d311, d214, d224);
	not (d312, d183);
	xor (d313, d221, d227);
	buf (d314, d125);
	buf (d315, d97);
	xnor (d316, d213, d231);
	or (d317, d224, d229);
	buf (d318, d74);
	and (d319, d218, d222);
	buf (d320, d186);
	nor (d321, d220, d228);
	nor (d322, d213, d220);
	not (d323, d184);
	xnor (d324, d215, d228);
	nor (d325, d214, d223);
	or (d326, d218, d225);
	buf (d327, d209);
	xnor (d328, d318, d320);
	buf (d329, d275);
	or (d330, d241, d314);
	xor (d331, d258, d278);
	xnor (d332, d253, d288);
	nand (d333, d303, d308);
	nor (d334, d260, d274);
	and (d335, d267, d321);
	or (d336, d304, d315);
	not (d337, d271);
	xor (d338, d269, d314);
	xor (d339, d238, d296);
	nor (d340, d239, d240);
	and (d341, d279, d295);
	buf (d342, d253);
	xor (d343, d273, d320);
	not (d344, d114);
	not (d345, d143);
	xnor (d346, d246, d306);
	nor (d347, d295, d303);
	nor (d348, d296, d320);
	nor (d349, d283, d293);
	or (d350, d241, d257);
	nand (d351, d304, d310);
	xor (d352, d311, d323);
	xnor (d353, d260, d269);
	not (d354, d310);
	and (d355, d273, d291);
	or (d356, d300, d318);
	xnor (d357, d250, d301);
	xnor (d358, d266, d306);
	not (d359, d182);
	and (d360, d244, d295);
	nor (d361, d247, d248);
	nand (d362, d312, d314);
	buf (d363, d181);
	xor (d364, d289, d305);
	not (d365, d49);
	not (d366, d110);
	not (d367, d127);
	xor (d368, d252, d273);
	xnor (d369, d241, d319);
	nor (d370, d297, d310);
	buf (d371, d304);
	not (d372, d28);
	not (d373, d98);
	not (d374, d219);
	xnor (d375, d283, d294);
	xor (d376, d246, d296);
	and (d377, d237, d316);
	xor (d378, d299, d308);
	nand (d379, d258, d296);
	xnor (d380, d272, d315);
	xor (d381, d273, d296);
	nand (d382, d278, d281);
	not (d383, d38);
	nor (d384, d278, d315);
	nor (d385, d264, d306);
	xnor (d386, d251, d256);
	or (d387, d309, d320);
	not (d388, d176);
	not (d389, d206);
	nor (d390, d275, d307);
	xnor (d391, d235, d271);
	and (d392, d284, d306);
	xnor (d393, d269, d304);
	xnor (d394, d249, d266);
	nor (d395, d255, d263);
	not (d396, d121);
	xnor (d397, d335, d344);
	or (d398, d351, d354);
	xnor (d399, d350, d392);
	buf (d400, d284);
	buf (d401, d383);
	and (d402, d389, d392);
	buf (d403, d212);
	xor (d404, d348);
	nand (d405, d340, d379);
	xor (d406, d347, d379);
	buf (d407, d135);
	buf (d408, d233);
	xor (d409, d341, d346);
	or (d410, d359, d364);
	not (d411, d329);
	and (d412, d328, d390);
	and (d413, d362, d392);
	nand (d414, d387, d393);
	and (d415, d337, d391);
	or (d416, d364, d367);
	and (d417, d337, d371);
	buf (d418, d98);
	and (d419, d336, d394);
	and (d420, d328, d341);
	buf (d421, d66);
	xor (d422, d402, d405);
	not (d423, d354);
	assign f1 = d422;
	assign f2 = d422;
	assign f3 = d422;
	assign f4 = d422;
	assign f5 = d422;
	assign f6 = d422;
	assign f7 = d422;
	assign f8 = d422;
endmodule
