module CCGRCG44( x0, x1, x2, x3, f1, f2, f3 );

	input x0, x1, x2, x3;
	output f1, f2, f3;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314, d315, d316, d317, d318, d319, d320, d321, d322, d323, d324, d325, d326, d327, d328, d329, d330, d331, d332, d333, d334, d335, d336, d337, d338, d339, d340, d341, d342, d343, d344, d345, d346, d347, d348, d349, d350, d351, d352, d353, d354, d355, d356, d357, d358, d359, d360, d361, d362, d363, d364, d365, d366, d367, d368, d369, d370, d371, d372, d373, d374, d375, d376, d377, d378, d379, d380, d381, d382, d383, d384, d385, d386, d387, d388, d389, d390, d391, d392, d393, d394, d395, d396, d397, d398, d399, d400, d401, d402, d403, d404, d405, d406, d407, d408, d409, d410, d411, d412, d413, d414, d415, d416, d417, d418, d419, d420, d421, d422, d423, d424, d425, d426, d427, d428, d429, d430, d431, d432, d433;

	nor (d1, x2, x3);
	nand (d2, x1);
	or (d3, x2, x3);
	or (d4, x0, x3);
	not (d5, x0);
	and (d6, x1, x2);
	or (d7, x1, x3);
	xnor (d8, x2, x3);
	xor (d9, x1);
	and (d10, x1, x3);
	xnor (d11, x0, x2);
	and (d12, x0);
	xor (d13, x1, x2);
	xnor (d14, x0, x2);
	or (d15, x2, x3);
	and (d16, x0, x1);
	not (d17, x3);
	and (d18, x2, x3);
	xnor (d19, x1, x3);
	nor (d20, x1, x2);
	or (d21, x1, x2);
	xor (d22, x0, x3);
	nand (d23, x0, x2);
	nor (d24, x2, x3);
	or (d25, x1, x2);
	buf (d26, x2);
	and (d27, x1);
	nor (d28, x1, x2);
	nor (d29, x0);
	xor (d30, x3);
	xor (d31, x0, x1);
	xor (d32, x0);
	nand (d33, x1, x3);
	xor (d34, x2, x3);
	nor (d35, x0, x1);
	nor (d36, x0, x2);
	nand (d37, x0);
	nand (d38, x0, x1);
	nand (d39, x0, x3);
	and (d40, x2);
	or (d41, d11, d14);
	or (d42, d15, d26);
	xnor (d43, d32, d39);
	or (d44, d4, d32);
	nor (d45, d8, d27);
	not (d46, d29);
	nand (d47, d31, d37);
	nand (d48, d2, d10);
	nor (d49, d9, d35);
	nand (d50, d20, d29);
	or (d51, d31, d33);
	buf (d52, d30);
	xor (d53, d31, d36);
	nand (d54, d5, d11);
	and (d55, d10, d24);
	xnor (d56, d1, d7);
	or (d57, d25, d36);
	nor (d58, d10, d34);
	xnor (d59, d29, d32);
	not (d60, d16);
	xor (d61, d13, d14);
	nor (d62, d17, d27);
	buf (d63, d24);
	and (d64, d8, d27);
	not (d65, d6);
	nor (d66, d14, d34);
	xor (d67, d5, d30);
	buf (d68, d25);
	not (d69, d61);
	buf (d70, d4);
	xor (d71, d50, d53);
	nand (d72, d59, d63);
	buf (d73, d29);
	and (d74, d61, d67);
	and (d75, d41, d67);
	and (d76, d41, d52);
	nand (d77, d45, d53);
	buf (d78, d41);
	not (d79, d47);
	xor (d80, d46, d58);
	xor (d81, d42, d45);
	not (d82, d55);
	xnor (d83, d47, d68);
	or (d84, d41, d46);
	nand (d85, d50, d65);
	xor (d86, d43, d62);
	buf (d87, d33);
	or (d88, d64, d67);
	buf (d89, d35);
	buf (d90, d51);
	buf (d91, d42);
	buf (d92, d31);
	nand (d93, d49, d68);
	xnor (d94, d44, d53);
	nor (d95, d43, d60);
	or (d96, d54, d61);
	buf (d97, d11);
	nor (d98, d42, d54);
	nand (d99, d41, d68);
	nand (d100, d45, d51);
	nor (d101, d57, d65);
	buf (d102, d13);
	nor (d103, d57, d59);
	xor (d104, d55, d63);
	and (d105, d54, d62);
	or (d106, d51, d56);
	not (d107, d30);
	and (d108, d44, d66);
	buf (d109, x3);
	xor (d110, d46, d49);
	or (d111, d65, d66);
	not (d112, d58);
	buf (d113, d12);
	or (d114, d56, d63);
	not (d115, d12);
	nand (d116, d45, d52);
	not (d117, d63);
	and (d118, d48, d63);
	or (d119, d57);
	and (d120, d43);
	nor (d121, d58, d59);
	or (d122, d67);
	and (d123, d52, d56);
	xnor (d124, d48, d58);
	xnor (d125, d54, d59);
	buf (d126, d68);
	or (d127, d52, d56);
	xnor (d128, d50, d51);
	nand (d129, d48, d64);
	or (d130, d41, d50);
	not (d131, d3);
	nand (d132, d47, d56);
	and (d133, d50, d54);
	not (d134, d13);
	nand (d135, d61, d68);
	xor (d136, d52, d57);
	not (d137, d10);
	xor (d138, d68);
	nand (d139, d46, d54);
	nor (d140, d46, d54);
	xnor (d141, d52, d65);
	nand (d142, d43, d56);
	xnor (d143, d62, d68);
	xor (d144, d41, d47);
	buf (d145, d59);
	xor (d146, d45, d47);
	nand (d147, d59, d64);
	xnor (d148, d74, d111);
	not (d149, d109);
	nor (d150, d74, d95);
	xor (d151, d82, d117);
	nor (d152, d86, d114);
	not (d153, d1);
	not (d154, d50);
	or (d155, d103, d108);
	nand (d156, d80, d125);
	not (d157, d134);
	xor (d158, d93, d113);
	xnor (d159, d84, d105);
	xor (d160, d78, d116);
	nand (d161, d72, d132);
	xnor (d162, d86, d117);
	not (d163, d22);
	xor (d164, d69, d104);
	xor (d165, d127, d139);
	or (d166, d104, d119);
	xnor (d167, d92, d125);
	and (d168, d102, d137);
	nor (d169, d94, d136);
	buf (d170, d134);
	and (d171, d71, d141);
	xor (d172, d98, d114);
	xnor (d173, d131, d136);
	nor (d174, d92, d136);
	buf (d175, d116);
	or (d176, d141, d145);
	xnor (d177, d85, d127);
	nor (d178, d70, d103);
	xnor (d179, d123, d126);
	not (d180, d65);
	xnor (d181, d87, d140);
	nand (d182, d158, d160);
	xor (d183, d157, d159);
	or (d184, d151, d176);
	nand (d185, d149, d171);
	not (d186, d54);
	not (d187, d66);
	xnor (d188, d172, d174);
	xnor (d189, d163, d175);
	xnor (d190, d166, d169);
	nand (d191, d150, d165);
	or (d192, d151, d152);
	and (d193, d165, d175);
	buf (d194, d104);
	and (d195, d161, d176);
	buf (d196, d90);
	nand (d197, d163, d165);
	not (d198, d155);
	or (d199, d150, d166);
	buf (d200, d117);
	and (d201, d151, d162);
	nor (d202, d159, d165);
	xnor (d203, d164, d172);
	xnor (d204, d148, d178);
	nor (d205, d155, d167);
	buf (d206, d84);
	nand (d207, d151, d158);
	xor (d208, d161, d178);
	nand (d209, d180, d181);
	xor (d210, d156, d161);
	nor (d211, d151, d179);
	not (d212, d52);
	not (d213, d108);
	xor (d214, d155, d173);
	nor (d215, d155, d162);
	xor (d216, d150, d173);
	or (d217, d152, d178);
	or (d218, d201, d206);
	buf (d219, d165);
	nor (d220, d198, d209);
	and (d221, d182, d202);
	nand (d222, d197, d215);
	nand (d223, d185, d196);
	xnor (d224, d185, d209);
	or (d225, d183, d213);
	buf (d226, d137);
	xor (d227, d202, d217);
	not (d228, d9);
	nand (d229, d186, d194);
	nor (d230, d195, d199);
	xor (d231, d182, d212);
	nor (d232, d183, d209);
	or (d233, d190, d196);
	and (d234, d186, d214);
	and (d235, d199, d210);
	nor (d236, d183, d188);
	not (d237, d143);
	nor (d238, d187, d199);
	or (d239, d202, d210);
	or (d240, d182, d210);
	xnor (d241, d182, d208);
	xor (d242, d211);
	or (d243, d189, d190);
	or (d244, d184, d212);
	nor (d245, d199, d214);
	nand (d246, d187, d192);
	and (d247, d209, d213);
	xor (d248, d196, d216);
	xor (d249, d191, d211);
	xor (d250, d190, d198);
	or (d251, d186, d198);
	or (d252, d185, d196);
	buf (d253, d154);
	or (d254, d188, d201);
	xor (d255, d186, d210);
	xnor (d256, d196, d206);
	xnor (d257, d199, d210);
	xor (d258, d191, d199);
	nor (d259, d196, d214);
	or (d260, d191, d193);
	nand (d261, d193, d210);
	xnor (d262, d189, d208);
	or (d263, d186, d194);
	and (d264, d195, d206);
	nor (d265, d199, d217);
	buf (d266, d48);
	nand (d267, d184, d214);
	xnor (d268, d189, d217);
	or (d269, d185, d186);
	nand (d270, d183, d193);
	not (d271, d110);
	not (d272, d36);
	and (d273, d189, d191);
	nand (d274, d186, d202);
	not (d275, d39);
	nand (d276, d202, d215);
	or (d277, d190, d217);
	not (d278, d112);
	nor (d279, d203, d206);
	and (d280, d185, d187);
	buf (d281, d53);
	or (d282, d200, d212);
	not (d283, d17);
	xnor (d284, d197, d199);
	not (d285, d32);
	xor (d286, d190, d204);
	nor (d287, d183, d212);
	or (d288, d190, d198);
	nor (d289, d213, d216);
	buf (d290, d179);
	nor (d291, d188, d213);
	or (d292, d182, d198);
	buf (d293, d45);
	xnor (d294, d205, d213);
	nand (d295, d193, d205);
	or (d296, d190, d207);
	nand (d297, d199, d203);
	xor (d298, d201, d210);
	xnor (d299, d206, d209);
	nor (d300, d196, d207);
	xnor (d301, d211, d217);
	or (d302, d237, d260);
	xor (d303, d255, d297);
	and (d304, d270, d299);
	nand (d305, d236, d237);
	not (d306, d221);
	xor (d307, d225, d290);
	or (d308, d221, d248);
	not (d309, d187);
	or (d310, d271, d288);
	or (d311, d218, d224);
	nand (d312, d247, d301);
	nor (d313, d248, d284);
	xor (d314, d277, d294);
	xnor (d315, d239, d283);
	xor (d316, d280, d284);
	nor (d317, d225, d298);
	buf (d318, d147);
	or (d319, d233, d265);
	xor (d320, d264, d293);
	nand (d321, d221, d236);
	and (d322, d263, d291);
	not (d323, d136);
	and (d324, d245, d292);
	not (d325, d106);
	xor (d326, d273, d280);
	nor (d327, d219, d300);
	nand (d328, d267, d288);
	or (d329, d259, d284);
	xor (d330, d223, d225);
	nor (d331, d246, d279);
	nand (d332, d271, d296);
	and (d333, d270, d272);
	buf (d334, d107);
	nor (d335, d246, d270);
	nand (d336, d226, d240);
	and (d337, d286, d297);
	xor (d338, d246, d258);
	xor (d339, d219, d267);
	nor (d340, d223, d300);
	xor (d341, d239, d279);
	not (d342, d277);
	or (d343, d259, d296);
	and (d344, d247, d274);
	not (d345, d201);
	nand (d346, d229, d239);
	nor (d347, d231, d243);
	xor (d348, d261, d267);
	nor (d349, d235, d272);
	or (d350, d226, d255);
	buf (d351, d62);
	xor (d352, d225, d297);
	or (d353, d244, d272);
	and (d354, d270, d295);
	not (d355, d177);
	and (d356, d266, d267);
	and (d357, d231, d260);
	nand (d358, d249, d259);
	not (d359, d86);
	buf (d360, d212);
	not (d361, d226);
	buf (d362, d230);
	xor (d363, d248, d268);
	buf (d364, d82);
	xor (d365, d254, d268);
	nand (d366, d231, d264);
	and (d367, d229, d280);
	nand (d368, d258, d272);
	nor (d369, d230, d253);
	buf (d370, d106);
	xor (d371, d230, d236);
	xor (d372, d219, d258);
	not (d373, d168);
	xor (d374, d246, d274);
	nand (d375, d282, d301);
	and (d376, d246, d267);
	nand (d377, d231, d238);
	xor (d378, d242, d263);
	not (d379, d252);
	nor (d380, d362);
	not (d381, d64);
	nor (d382, d362, d363);
	and (d383, d334, d338);
	and (d384, d360, d373);
	and (d385, d335, d354);
	nand (d386, d332, d344);
	nor (d387, d331, d341);
	xnor (d388, d348, d366);
	and (d389, d309, d370);
	xnor (d390, d340, d375);
	buf (d391, d49);
	nor (d392, d317, d379);
	and (d393, d349, d355);
	nand (d394, d334, d340);
	nor (d395, d336, d350);
	nand (d396, d353, d365);
	not (d397, d369);
	or (d398, d354, d355);
	xnor (d399, d305, d310);
	or (d400, d329, d377);
	nor (d401, d330, d334);
	xnor (d402, d314, d338);
	nand (d403, d311, d370);
	or (d404, d317, d351);
	and (d405, d353, d360);
	nor (d406, d341, d370);
	or (d407, d319, d339);
	nor (d408, d329, d350);
	or (d409, d323, d352);
	and (d410, d356, d375);
	nor (d411, d307, d341);
	xnor (d412, d361, d369);
	nor (d413, d312, d360);
	or (d414, d315, d319);
	nor (d415, d306, d329);
	nand (d416, d355, d370);
	xnor (d417, d307, d316);
	and (d418, d320, d353);
	or (d419, d308, d350);
	and (d420, d332, d356);
	nor (d421, d309, d352);
	and (d422, d348, d356);
	buf (d423, d327);
	or (d424, d339, d350);
	buf (d425, d274);
	nor (d426, d332, d378);
	and (d427, d346, d367);
	xor (d428, d323, d356);
	or (d429, d308, d338);
	and (d430, d305, d340);
	buf (d431, d284);
	or (d432, d304, d374);
	nand (d433, d302, d315);
	assign f1 = d432;
	assign f2 = d420;
	assign f3 = d402;
endmodule
