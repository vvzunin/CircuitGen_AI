module CCGRCG184( x0, x1, x2, x3, x4, x5, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17, f18 );

	input x0, x1, x2, x3, x4, x5;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17, f18;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314, d315, d316, d317, d318, d319, d320, d321, d322, d323, d324, d325, d326, d327, d328, d329, d330, d331, d332, d333, d334, d335, d336, d337, d338, d339, d340, d341, d342, d343, d344, d345, d346, d347, d348, d349, d350, d351, d352, d353, d354, d355, d356, d357, d358, d359, d360, d361, d362, d363, d364, d365, d366, d367, d368, d369, d370, d371, d372, d373, d374, d375, d376, d377, d378, d379, d380, d381, d382, d383, d384, d385, d386, d387, d388, d389, d390, d391, d392, d393, d394, d395;

	not (d1, x1);
	and (d2, x0);
	nor (d3, x0, x3);
	buf (d4, x5);
	and (d5, x1, x2);
	nand (d6, x3, x4);
	xor (d7, x2, x5);
	xor (d8, x1, x5);
	nand (d9, x2, x3);
	and (d10, x2, x5);
	xnor (d11, x0, x5);
	buf (d12, x0);
	buf (d13, x2);
	and (d14, x5);
	nor (d15, x3);
	xnor (d16, x5);
	not (d17, x2);
	xnor (d18, x0, x2);
	buf (d19, x4);
	and (d20, x0, x3);
	xnor (d21, x0, x3);
	and (d22, x3, x5);
	xnor (d23, x2, x5);
	xor (d24, x1, x3);
	and (d25, x1, x5);
	or (d26, x0, x3);
	xnor (d27, x4, x5);
	not (d28, x5);
	xnor (d29, x3, x4);
	nor (d30, x5);
	and (d31, x0, x2);
	and (d32, x1, x4);
	and (d33, x4);
	xor (d34, x2, x3);
	nand (d35, x0, x5);
	or (d36, x1, x4);
	or (d37, x0, x1);
	xnor (d38, x1, x2);
	buf (d39, x3);
	xor (d40, x1, x4);
	or (d41, x1, x2);
	nor (d42, x4, x5);
	or (d43, x1, x3);
	xor (d44, x0, x2);
	xor (d45, x0, x1);
	xor (d46, x2, x4);
	not (d47, x0);
	xor (d48, x2, x5);
	nand (d49, x2);
	and (d50, x3);
	or (d51, x2);
	or (d52, x2, x4);
	nand (d53, x4, x5);
	and (d54, x3, x4);
	or (d55, x4);
	xnor (d56, x0, x4);
	xnor (d57, x1, x3);
	not (d58, d18);
	nor (d59, d16, d23);
	not (d60, d9);
	buf (d61, d52);
	buf (d62, d39);
	nor (d63, d32, d53);
	not (d64, x4);
	nand (d65, d27, d33);
	and (d66, d11, d44);
	nand (d67, d5, d24);
	and (d68, d13, d33);
	not (d69, d48);
	not (d70, d19);
	xnor (d71, d47, d48);
	nor (d72, d5, d30);
	buf (d73, d45);
	xnor (d74, d12, d25);
	nand (d75, d31, d53);
	nand (d76, d18, d33);
	xnor (d77, d23, d36);
	and (d78, d36, d40);
	xor (d79, d3, d35);
	and (d80, d5, d55);
	xor (d81, d6, d56);
	xnor (d82, d24, d31);
	nand (d83, d10, d38);
	xor (d84, d22, d43);
	not (d85, d17);
	and (d86, d5, d11);
	or (d87, d30, d42);
	nand (d88, d24, d42);
	not (d89, d28);
	nand (d90, d36, d43);
	buf (d91, d34);
	buf (d92, d56);
	xor (d93, d38, d47);
	not (d94, d36);
	or (d95, d30, d51);
	nor (d96, d8, d11);
	xor (d97, d41, d54);
	xor (d98, d20, d45);
	buf (d99, d22);
	nand (d100, d45, d57);
	or (d101, d14, d45);
	xnor (d102, d20, d22);
	xor (d103, d37, d55);
	or (d104, d3, d41);
	nand (d105, d4, d17);
	and (d106, d47, d55);
	xor (d107, d39, d44);
	xnor (d108, d31, d46);
	nand (d109, d9, d22);
	nor (d110, d22, d51);
	and (d111, d79, d98);
	xnor (d112, d81, d109);
	nor (d113, d88, d93);
	not (d114, d27);
	xnor (d115, d101, d110);
	buf (d116, d64);
	nor (d117, d75, d93);
	and (d118, d73, d76);
	not (d119, d81);
	nor (d120, d68, d81);
	nor (d121, d69, d108);
	not (d122, d63);
	nand (d123, d67, d100);
	xor (d124, d62, d86);
	buf (d125, d21);
	and (d126, d79, d92);
	xnor (d127, d84, d85);
	and (d128, d70, d106);
	xor (d129, d97, d98);
	nor (d130, d61, d85);
	and (d131, d77, d104);
	or (d132, d84, d103);
	buf (d133, d32);
	xnor (d134, d95, d107);
	not (d135, d10);
	xor (d136, d71, d107);
	or (d137, d83, d91);
	not (d138, d72);
	or (d139, d67, d69);
	not (d140, d107);
	nor (d141, d81, d85);
	and (d142, d77, d94);
	or (d143, d76, d102);
	xnor (d144, d87, d91);
	or (d145, d77, d88);
	xor (d146, d62, d86);
	nor (d147, d58, d81);
	buf (d148, d74);
	buf (d149, d68);
	not (d150, d90);
	or (d151, d66, d72);
	xnor (d152, d66, d101);
	nand (d153, d86, d90);
	nand (d154, d81, d94);
	buf (d155, d46);
	or (d156, d80, d91);
	not (d157, d31);
	xor (d158, d99, d103);
	buf (d159, d55);
	xnor (d160, d144, d146);
	and (d161, d114, d131);
	nor (d162, d123, d143);
	xnor (d163, d112, d134);
	xnor (d164, d126, d144);
	or (d165, d140, d153);
	buf (d166, d66);
	and (d167, d141, d151);
	xor (d168, d139, d157);
	nor (d169, d142, d158);
	nand (d170, d113, d135);
	and (d171, d130, d131);
	nand (d172, d119, d120);
	or (d173, d145, d150);
	xnor (d174, d131, d132);
	xnor (d175, d123, d142);
	nor (d176, d132, d138);
	nor (d177, d124, d149);
	nand (d178, d124, d148);
	or (d179, d124, d139);
	and (d180, d122, d144);
	xnor (d181, d113, d120);
	nand (d182, d120, d140);
	nor (d183, d149, d155);
	xor (d184, d155, d156);
	buf (d185, d150);
	and (d186, d131, d157);
	xor (d187, d135, d142);
	xor (d188, d117, d134);
	buf (d189, d12);
	buf (d190, d26);
	xnor (d191, d130, d141);
	nand (d192, d134, d146);
	nor (d193, d127, d141);
	nand (d194, d131, d143);
	and (d195, d153, d155);
	xnor (d196, d135, d151);
	xnor (d197, d118, d155);
	nand (d198, d133, d138);
	buf (d199, d146);
	and (d200, d118, d120);
	nand (d201, d128, d154);
	xor (d202, d135, d154);
	nand (d203, d120, d148);
	buf (d204, d125);
	xor (d205, d111, d113);
	nor (d206, d116, d154);
	or (d207, d131, d157);
	xnor (d208, d143, d154);
	nand (d209, d140, d145);
	and (d210, d118, d158);
	and (d211, d143, d156);
	nor (d212, d127, d140);
	nor (d213, d124, d138);
	not (d214, d51);
	buf (d215, d44);
	and (d216, d121, d152);
	nand (d217, d140, d157);
	nand (d218, d139, d156);
	xor (d219, d113, d131);
	buf (d220, d71);
	nor (d221, d137, d154);
	nor (d222, d127, d149);
	or (d223, d124, d138);
	xnor (d224, d116, d129);
	and (d225, d130, d152);
	xnor (d226, d154);
	and (d227, d112, d143);
	xor (d228, d112, d121);
	nand (d229, d123, d141);
	nand (d230, d154, d155);
	or (d231, d147, d150);
	or (d232, d136, d138);
	xnor (d233, d125, d153);
	xnor (d234, d147, d154);
	xnor (d235, d129, d156);
	xnor (d236, d118, d123);
	not (d237, d91);
	nor (d238, d136);
	buf (d239, d17);
	nor (d240, d139, d148);
	nand (d241, d131, d154);
	not (d242, d35);
	nor (d243, d122, d123);
	buf (d244, d234);
	nor (d245, d217, d236);
	xor (d246, d193, d240);
	buf (d247, d51);
	nor (d248, d178, d194);
	and (d249, d173, d208);
	and (d250, d189);
	xnor (d251, d196, d219);
	nand (d252, d194, d215);
	nand (d253, d171, d190);
	xnor (d254, d164, d213);
	not (d255, d69);
	and (d256, d190, d192);
	not (d257, d155);
	not (d258, d23);
	xor (d259, d174, d190);
	nor (d260, d194, d228);
	buf (d261, d149);
	xor (d262, d175, d215);
	buf (d263, d58);
	xnor (d264, d189, d223);
	buf (d265, d89);
	and (d266, d179, d222);
	nor (d267, d164, d225);
	or (d268, d186, d192);
	xnor (d269, d177, d243);
	nor (d270, d262, d266);
	not (d271, d15);
	nand (d272, d245, d250);
	xnor (d273, d252, d267);
	xor (d274, d260, d261);
	buf (d275, d30);
	or (d276, d270, d274);
	nor (d277, d272);
	xnor (d278, d270, d272);
	buf (d279, d73);
	buf (d280, d119);
	buf (d281, d141);
	and (d282, d271, d274);
	nand (d283, d272, d274);
	or (d284, d272);
	not (d285, d25);
	nand (d286, d270, d271);
	or (d287, d270, d271);
	xor (d288, d271, d273);
	nand (d289, d273, d274);
	nor (d290, d270, d272);
	not (d291, d57);
	or (d292, d270, d272);
	and (d293, d270, d273);
	buf (d294, d49);
	xnor (d295, d274);
	nand (d296, d270, d271);
	and (d297, d270, d272);
	xor (d298, d270, d274);
	xnor (d299, d272, d273);
	and (d300, d274);
	nor (d301, d271);
	xnor (d302, d272, d274);
	nor (d303, d270, d272);
	or (d304, d270, d271);
	and (d305, d272, d274);
	nand (d306, d270, d274);
	buf (d307, d200);
	not (d308, d8);
	xor (d309, d271);
	nand (d310, d271, d272);
	nor (d311, d271, d274);
	buf (d312, d158);
	nor (d313, d271, d273);
	nand (d314, d270, d273);
	nor (d315, d270, d274);
	nor (d316, d273);
	buf (d317, d133);
	nand (d318, d272, d273);
	or (d319, d272, d274);
	xor (d320, d274);
	or (d321, d271, d274);
	or (d322, d271);
	nor (d323, d270, d273);
	or (d324, d273, d274);
	buf (d325, d69);
	xor (d326, d270, d273);
	and (d327, d270, d274);
	or (d328, d302, d316);
	xnor (d329, d298, d299);
	or (d330, d298, d312);
	not (d331, d29);
	xor (d332, d303, d326);
	xnor (d333, d284, d327);
	xnor (d334, d318, d319);
	xnor (d335, d314, d320);
	nor (d336, d318, d326);
	xor (d337, d311, d314);
	xor (d338, d276, d310);
	not (d339, d93);
	buf (d340, d317);
	not (d341, d243);
	and (d342, d306, d311);
	and (d343, d284, d312);
	or (d344, d293, d303);
	nor (d345, d293, d322);
	or (d346, d326);
	and (d347, d275, d316);
	nor (d348, d278, d327);
	buf (d349, d318);
	nand (d350, d331, d346);
	nor (d351, d334, d339);
	xor (d352, d332, d345);
	not (d353, d30);
	buf (d354, d148);
	not (d355, d89);
	and (d356, d342, d349);
	xor (d357, d339, d347);
	xor (d358, d337, d346);
	not (d359, d313);
	not (d360, d219);
	not (d361, d130);
	nand (d362, d331, d334);
	and (d363, d331, d332);
	not (d364, d189);
	buf (d365, d109);
	xor (d366, d341, d349);
	xor (d367, d331, d332);
	not (d368, d182);
	xnor (d369, d336, d342);
	or (d370, d331, d346);
	and (d371, d344);
	or (d372, d338, d349);
	nor (d373, d337, d346);
	or (d374, d335, d347);
	or (d375, d331, d343);
	nand (d376, d330, d332);
	not (d377, d304);
	not (d378, d98);
	and (d379, d329, d334);
	and (d380, d330, d332);
	and (d381, d328, d331);
	xor (d382, d344, d347);
	nor (d383, d330, d336);
	xor (d384, d340, d346);
	nor (d385, d336, d342);
	nor (d386, d333, d346);
	or (d387, d328, d346);
	nand (d388, d332, d348);
	not (d389, d172);
	or (d390, d332, d337);
	or (d391, d331, d333);
	nor (d392, d341, d347);
	nand (d393, d337, d342);
	buf (d394, d181);
	and (d395, d331, d334);
	assign f1 = d390;
	assign f2 = d376;
	assign f3 = d372;
	assign f4 = d374;
	assign f5 = d352;
	assign f6 = d354;
	assign f7 = d379;
	assign f8 = d358;
	assign f9 = d381;
	assign f10 = d379;
	assign f11 = d373;
	assign f12 = d393;
	assign f13 = d366;
	assign f14 = d394;
	assign f15 = d350;
	assign f16 = d389;
	assign f17 = d366;
	assign f18 = d384;
endmodule
