module CCGRCG181( x0, x1, x2, x3, x4, x5, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16 );

	input x0, x1, x2, x3, x4, x5;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314, d315, d316, d317, d318, d319, d320, d321, d322, d323, d324, d325, d326, d327, d328, d329, d330;

	or (d1, x0, x3);
	and (d2, x2, x5);
	nor (d3, x1, x4);
	nor (d4, x1, x2);
	and (d5, x0, x2);
	buf (d6, x1);
	and (d7, x0, x5);
	nand (d8, x1, x2);
	nor (d9, x0, x2);
	or (d10, x0, x3);
	nor (d11, x3, x4);
	buf (d12, x0);
	xor (d13, x0, x2);
	or (d14, x2, x3);
	xor (d15, x0, x1);
	or (d16, x3, x5);
	nand (d17, x0, x1);
	and (d18, x3, x5);
	xor (d19, x2);
	not (d20, x5);
	xor (d21, x1, x3);
	xor (d22, x5);
	or (d23, x0, x1);
	nand (d24, x5);
	xnor (d25, x1, x2);
	or (d26, x1, x3);
	or (d27, x5);
	not (d28, x3);
	nand (d29, x4);
	buf (d30, x3);
	xnor (d31, x0, x2);
	nand (d32, x1);
	and (d33, x3, x4);
	nor (d34, x2, x3);
	nand (d35, x2);
	and (d36, x1, x4);
	not (d37, x1);
	or (d38, x0, x4);
	and (d39, x1, x5);
	or (d40, x1, x5);
	xor (d41, x1, x4);
	nand (d42, x3, x4);
	buf (d43, x4);
	and (d44, x4);
	buf (d45, x5);
	and (d46, x3, x4);
	xor (d47, x1, x3);
	xnor (d48, x2, x4);
	xor (d49, x0, x3);
	xnor (d50, x4, x5);
	nor (d51, x2, x4);
	buf (d52, x2);
	not (d53, x4);
	nor (d54, x0, x1);
	and (d55, x0, x3);
	nand (d56, x0, x3);
	xor (d57, x0, x5);
	not (d58, d5);
	or (d59, d5, d35);
	xnor (d60, d24, d48);
	nor (d61, d29, d57);
	not (d62, d7);
	and (d63, d29, d51);
	buf (d64, d4);
	nand (d65, d13, d14);
	buf (d66, d32);
	nor (d67, d11, d41);
	nand (d68, d14, d46);
	xnor (d69, d16);
	and (d70, d22);
	nor (d71, d37, d42);
	not (d72, d37);
	and (d73, d11, d40);
	xor (d74, d11, d35);
	nor (d75, d42, d49);
	nor (d76, d11, d22);
	and (d77, d26, d49);
	or (d78, d32, d33);
	or (d79, d10, d23);
	nor (d80, d10, d34);
	buf (d81, d2);
	xnor (d82, d22, d24);
	and (d83, d5, d49);
	not (d84, d39);
	nand (d85, d27, d41);
	and (d86, d18, d22);
	not (d87, d42);
	buf (d88, d28);
	xnor (d89, d31, d39);
	xor (d90, d19, d40);
	and (d91, d9, d31);
	or (d92, d11, d24);
	nor (d93, d15, d36);
	buf (d94, d52);
	nor (d95, d13, d53);
	nor (d96, d1, d29);
	xor (d97, d26, d39);
	or (d98, d49, d52);
	or (d99, d26, d37);
	xor (d100, d29, d52);
	buf (d101, d27);
	or (d102, d36, d47);
	or (d103, d13, d53);
	and (d104, d4, d31);
	nor (d105, d12, d44);
	xnor (d106, d38, d55);
	not (d107, d1);
	nand (d108, d16, d45);
	nand (d109, d5, d55);
	buf (d110, d46);
	xnor (d111, d31, d49);
	nor (d112, d20, d30);
	buf (d113, d54);
	not (d114, d51);
	xor (d115, d28, d33);
	not (d116, d11);
	buf (d117, d47);
	and (d118, d44, d46);
	and (d119, d4, d9);
	not (d120, d49);
	xnor (d121, d4, d5);
	xnor (d122, d21, d43);
	or (d123, d7, d54);
	or (d124, d20, d55);
	xor (d125, d41, d48);
	and (d126, d5, d49);
	buf (d127, d16);
	xor (d128, d10, d54);
	xnor (d129, d12, d16);
	xnor (d130, d11, d45);
	or (d131, d20, d35);
	nand (d132, d33, d41);
	nor (d133, d4, d45);
	not (d134, d16);
	nor (d135, d39, d51);
	buf (d136, d37);
	and (d137, d48, d49);
	xor (d138, d4, d20);
	xnor (d139, d12, d21);
	xnor (d140, d34, d56);
	buf (d141, d25);
	nor (d142, d11, d53);
	buf (d143, d34);
	nand (d144, d94, d120);
	nor (d145, d77, d123);
	nand (d146, d96, d138);
	xnor (d147, d59, d140);
	not (d148, d99);
	xor (d149, d132, d133);
	not (d150, d4);
	buf (d151, d6);
	not (d152, d96);
	buf (d153, d39);
	or (d154, d82, d92);
	nand (d155, d76, d87);
	nand (d156, d120, d125);
	xor (d157, d113, d137);
	xnor (d158, d119, d127);
	not (d159, d31);
	xnor (d160, d58, d89);
	nor (d161, d70, d92);
	xnor (d162, d80, d90);
	nand (d163, d136, d137);
	not (d164, d9);
	xor (d165, d58, d60);
	or (d166, d99, d128);
	nand (d167, d81, d90);
	nand (d168, d126, d137);
	xnor (d169, d61, d134);
	xnor (d170, d157, d168);
	nand (d171, d148, d157);
	xor (d172, d147, d164);
	xor (d173, d155, d160);
	xor (d174, d150, d167);
	nor (d175, d154, d158);
	not (d176, d22);
	nor (d177, d145, d159);
	buf (d178, d21);
	xor (d179, d156, d158);
	nor (d180, d151, d154);
	xnor (d181, d150, d152);
	buf (d182, d95);
	xor (d183, d158, d160);
	nor (d184, d159, d166);
	xor (d185, d148, d151);
	not (d186, d13);
	and (d187, d158, d163);
	xnor (d188, d143, d154);
	or (d189, d149, d160);
	not (d190, d169);
	or (d191, d150, d152);
	nor (d192, d146, d150);
	nor (d193, d160);
	and (d194, d148, d150);
	nor (d195, d156, d162);
	nand (d196, d146, d164);
	or (d197, d154, d165);
	buf (d198, d29);
	buf (d199, d44);
	nand (d200, d153, d162);
	xor (d201, d149, d154);
	xor (d202, d148);
	nand (d203, d146, d155);
	xnor (d204, d143, d148);
	nor (d205, d146, d161);
	or (d206, d162, d164);
	or (d207, d157, d165);
	nand (d208, d145, d166);
	nand (d209, d148, d168);
	nor (d210, d144, d148);
	or (d211, d164, d168);
	nor (d212, d148, d165);
	xnor (d213, d143, d164);
	nand (d214, d147, d160);
	nor (d215, d167, d169);
	nand (d216, d156, d169);
	or (d217, d151, d155);
	or (d218, d143, d153);
	xnor (d219, d161, d162);
	nor (d220, d144, d161);
	xnor (d221, d159, d164);
	xor (d222, d143, d148);
	nand (d223, d151, d162);
	xor (d224, d149, d150);
	nor (d225, d145, d160);
	nand (d226, d143, d154);
	and (d227, d145, d160);
	or (d228, d154, d161);
	not (d229, d78);
	nand (d230, d145, d165);
	xnor (d231, d148, d169);
	and (d232, d152, d155);
	nor (d233, d150, d166);
	and (d234, d148, d166);
	buf (d235, d69);
	or (d236, d156, d165);
	not (d237, d153);
	or (d238, d174, d200);
	or (d239, d176, d230);
	xor (d240, d185, d233);
	xor (d241, d180, d225);
	nand (d242, d174, d232);
	and (d243, d222, d234);
	and (d244, d200, d226);
	xnor (d245, d171, d181);
	xnor (d246, d185, d224);
	nand (d247, d188, d211);
	nand (d248, d212, d222);
	nor (d249, d178, d189);
	or (d250, d172, d199);
	nand (d251, d206, d231);
	not (d252, d150);
	xor (d253, d237, d251);
	xnor (d254, d245, d250);
	xor (d255, d250, d251);
	and (d256, d240, d242);
	nor (d257, d244, d251);
	not (d258, d208);
	xor (d259, d237, d241);
	not (d260, d116);
	and (d261, d238, d241);
	buf (d262, d111);
	nor (d263, d241, d242);
	not (d264, d20);
	nand (d265, d239, d251);
	xor (d266, d242, d246);
	buf (d267, d17);
	or (d268, d243, d250);
	nand (d269, d239, d245);
	nand (d270, d243, d246);
	or (d271, d237, d251);
	nor (d272, d247, d248);
	xor (d273, d237, d238);
	nor (d274, d243, d247);
	not (d275, d25);
	nor (d276, d237, d244);
	buf (d277, d10);
	not (d278, d94);
	or (d279, d240, d244);
	nor (d280, d239, d246);
	buf (d281, d124);
	nor (d282, d245, d249);
	nand (d283, d239, d242);
	or (d284, d242, d243);
	nor (d285, d267, d275);
	nand (d286, d256, d275);
	or (d287, d261, d284);
	buf (d288, d247);
	nand (d289, d286, d287);
	not (d290, d227);
	nor (d291, d285, d286);
	and (d292, d285, d287);
	or (d293, d285, d287);
	buf (d294, d224);
	nand (d295, d286, d287);
	xor (d296, d287, d288);
	xnor (d297, d287, d288);
	nand (d298, d286, d288);
	and (d299, d285, d288);
	and (d300, d286, d288);
	nor (d301, d287);
	nor (d302, d285);
	not (d303, d225);
	or (d304, d285, d287);
	or (d305, d286);
	not (d306, d170);
	nand (d307, d287, d288);
	and (d308, d285, d287);
	or (d309, d285, d286);
	or (d310, d286, d287);
	and (d311, d286, d287);
	or (d312, d285, d286);
	buf (d313, d274);
	and (d314, d285, d288);
	not (d315, d223);
	buf (d316, d179);
	and (d317, d286, d288);
	and (d318, d286);
	xor (d319, d286, d288);
	xnor (d320, d285, d286);
	buf (d321, d107);
	and (d322, d287, d288);
	nor (d323, d285, d288);
	buf (d324, d94);
	not (d325, d217);
	or (d326, d285, d288);
	nand (d327, d286, d288);
	and (d328, d287, d288);
	xor (d329, d286, d287);
	or (d330, d287);
	assign f1 = d289;
	assign f2 = d295;
	assign f3 = d325;
	assign f4 = d307;
	assign f5 = d299;
	assign f6 = d299;
	assign f7 = d303;
	assign f8 = d325;
	assign f9 = d296;
	assign f10 = d307;
	assign f11 = d304;
	assign f12 = d315;
	assign f13 = d320;
	assign f14 = d300;
	assign f15 = d298;
	assign f16 = d328;
endmodule
