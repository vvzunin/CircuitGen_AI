module CCGRCG51( x0, x1, x2, f1, f2, f3, f4, f5, f6, f7, f8 );

	input x0, x1, x2;
	output f1, f2, f3, f4, f5, f6, f7, f8;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104;

	nor (d1, x0, x1);
	and (d2, x1, x2);
	not (d3, x0);
	nand (d4, x0, x2);
	nand (d5, x1, x2);
	or (d6, x2);
	nand (d7, x1);
	xnor (d8, x1, x2);
	nor (d9, x1, x2);
	nor (d10, x1, x2);
	or (d11, x0, x2);
	xor (d12, x2);
	xor (d13, x0, x1);
	buf (d14, x1);
	or (d15, x1);
	xnor (d16, x0, x1);
	and (d17, x0, x2);
	nand (d18, x1, x2);
	xnor (d19, x1, x2);
	xnor (d20, x2);
	xnor (d21, x0, x1);
	nor (d22, x0, x2);
	nand (d23, x0, x1);
	xor (d24, x1, x2);
	not (d25, x1);
	and (d26, x0, x1);
	nor (d27, x1);
	xor (d28, x1);
	not (d29, x2);
	buf (d30, x0);
	nor (d31, x2);
	and (d32, x0);
	nand (d33, x0);
	nor (d34, x0, x1);
	and (d35, x0, x2);
	or (d36, x1, x2);
	and (d37, x1, x2);
	nor (d38, x0);
	xnor (d39, x1);
	xnor (d40, x0, x2);
	buf (d41, x2);
	not (d42, d12);
	xnor (d43, d18, d36);
	xor (d44, d3, d16);
	buf (d45, d36);
	buf (d46, d28);
	xor (d47, d15, d27);
	nor (d48, d19, d41);
	nand (d49, d28, d29);
	buf (d50, d1);
	nor (d51, d2, d33);
	not (d52, d41);
	buf (d53, d2);
	xnor (d54, d35, d41);
	xor (d55, d6, d23);
	nor (d56, d12, d19);
	nand (d57, d10, d17);
	or (d58, d37, d39);
	not (d59, d38);
	not (d60, d19);
	buf (d61, d21);
	not (d62, d26);
	nand (d63, d17, d28);
	or (d64, d3, d7);
	or (d65, d16);
	nor (d66, d16, d34);
	and (d67, d17, d21);
	buf (d68, d3);
	xor (d69, d23, d27);
	or (d70, d6, d15);
	xor (d71, d8, d15);
	xor (d72, d11, d31);
	nand (d73, d4, d39);
	not (d74, d28);
	or (d75, d15, d41);
	and (d76, d29, d32);
	xnor (d77, d3, d8);
	nand (d78, d28, d37);
	not (d79, d39);
	buf (d80, d34);
	xnor (d81, d15, d35);
	buf (d82, d14);
	nor (d83, d1, d25);
	buf (d84, d5);
	and (d85, d26);
	xor (d86, d17, d19);
	xnor (d87, d7, d25);
	not (d88, d33);
	nand (d89, d30, d36);
	xor (d90, d11, d24);
	nor (d91, d5, d27);
	or (d92, d13, d22);
	nand (d93, d9, d16);
	nand (d94, d11, d38);
	nand (d95, d35, d40);
	and (d96, d28, d41);
	buf (d97, d22);
	nand (d98, d26, d33);
	or (d99, d19, d24);
	or (d100, d7, d30);
	xnor (d101, d22, d30);
	and (d102, d12, d23);
	and (d103, d2, d8);
	xnor (d104, d6, d24);
	assign f1 = d63;
	assign f2 = d73;
	assign f3 = d47;
	assign f4 = d95;
	assign f5 = d55;
	assign f6 = d96;
	assign f7 = d101;
	assign f8 = d73;
endmodule
