module CCGRCG129( x0, x1, x2, x3, x4, f1, f2, f3, f4, f5, f6, f7, f8, f9 );

	input x0, x1, x2, x3, x4;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314, d315, d316, d317, d318, d319, d320, d321, d322, d323, d324, d325, d326, d327, d328, d329, d330, d331, d332, d333, d334, d335, d336, d337, d338, d339, d340, d341, d342, d343, d344, d345, d346, d347, d348, d349, d350, d351, d352, d353, d354, d355, d356, d357, d358, d359, d360, d361, d362, d363, d364, d365, d366, d367, d368, d369, d370, d371, d372, d373, d374, d375, d376, d377, d378, d379, d380, d381, d382, d383, d384, d385, d386, d387, d388, d389, d390, d391, d392, d393, d394, d395, d396, d397, d398, d399, d400, d401, d402, d403, d404, d405, d406, d407, d408, d409, d410, d411, d412, d413, d414, d415, d416, d417, d418, d419, d420, d421, d422, d423, d424, d425, d426, d427, d428, d429, d430, d431, d432, d433, d434, d435, d436, d437, d438, d439, d440, d441, d442, d443, d444, d445, d446, d447, d448, d449, d450, d451, d452, d453, d454, d455, d456, d457, d458, d459, d460, d461, d462, d463, d464, d465, d466, d467, d468, d469, d470, d471, d472, d473, d474, d475, d476, d477, d478, d479, d480, d481, d482, d483, d484, d485, d486, d487, d488, d489, d490, d491, d492, d493, d494, d495;

	xor (d1, x4);
	nand (d2, x1);
	not (d3, x4);
	and (d4, x0, x2);
	buf (d5, x0);
	nand (d6, x2);
	and (d7, x1, x3);
	not (d8, x2);
	and (d9, x3, x4);
	nor (d10, x0, x2);
	or (d11, x0, x1);
	xnor (d12, x0, x2);
	or (d13, x1, x2);
	buf (d14, x2);
	xor (d15, x0, x4);
	and (d16, x2);
	and (d17, x0);
	or (d18, x0, x3);
	xor (d19, x1, x3);
	or (d20, x4);
	xnor (d21, x1, x2);
	xor (d22, x2, x4);
	nor (d23, x0, x4);
	buf (d24, x3);
	buf (d25, x1);
	xnor (d26, x2, x3);
	nor (d27, x1, x3);
	or (d28, x0, x2);
	nor (d29, x0, x1);
	xnor (d30, x0, x4);
	not (d31, x1);
	nand (d32, x0, x4);
	or (d33, x2, x4);
	and (d34, x0, x3);
	xor (d35, x0, x3);
	nand (d36, x0, x3);
	nor (d37, x1, x4);
	nor (d38, x2, x3);
	nand (d39, x0, x4);
	nand (d40, x0, x3);
	xor (d41, x1, x2);
	nor (d42, x0);
	or (d43, x3, x4);
	or (d44, x0, x2);
	or (d45, x1, x3);
	nand (d46, x3);
	not (d47, x3);
	nor (d48, x3, x4);
	xor (d49, x0, x2);
	nand (d50, x0);
	and (d51, x2, x4);
	or (d52, x2);
	xor (d53, x0);
	xor (d54, x2, x4);
	nand (d55, x2, x3);
	and (d56, x2, x3);
	xnor (d57, x0, x3);
	nor (d58, x2, x4);
	buf (d59, x4);
	nor (d60, x0, x1);
	and (d61, x0, x2);
	nor (d62, x3, x4);
	xnor (d63, x0, x1);
	or (d64, x2, x4);
	xnor (d65, x2, x4);
	buf (d66, d35);
	not (d67, d52);
	and (d68, d33, d44);
	buf (d69, d28);
	or (d70, d22, d64);
	nor (d71, d9, d20);
	buf (d72, d19);
	or (d73, d45, d53);
	or (d74, d23, d53);
	nand (d75, d7, d58);
	nor (d76, d25, d39);
	xor (d77, d2, d5);
	nand (d78, d32, d53);
	nor (d79, d25, d58);
	nor (d80, d26, d56);
	nand (d81, d59);
	nor (d82, d11, d60);
	buf (d83, d34);
	xnor (d84, d8, d63);
	and (d85, d29, d64);
	nor (d86, d13, d32);
	and (d87, d29, d63);
	nand (d88, d23, d28);
	xnor (d89, d39, d50);
	nor (d90, d10, d28);
	or (d91, d16, d30);
	nand (d92, d74, d79);
	buf (d93, d42);
	xor (d94, d71, d76);
	and (d95, d68, d78);
	or (d96, d74, d84);
	nand (d97, d68, d90);
	or (d98, d70, d74);
	nor (d99, d67, d68);
	not (d100, d49);
	nand (d101, d68, d77);
	nand (d102, d66, d81);
	and (d103, d69, d71);
	nand (d104, d81, d91);
	nand (d105, d78, d86);
	xor (d106, d72, d87);
	and (d107, d76, d83);
	nor (d108, d69, d79);
	nor (d109, d71, d89);
	xor (d110, d72, d89);
	nor (d111, d77, d88);
	nor (d112, d67, d84);
	or (d113, d68, d84);
	nand (d114, d67, d84);
	xor (d115, d79, d84);
	nand (d116, d76, d91);
	nand (d117, d68, d91);
	not (d118, d10);
	xnor (d119, d77, d82);
	nor (d120, d69, d75);
	xor (d121, d74, d86);
	not (d122, d63);
	xor (d123, d72, d88);
	buf (d124, d48);
	xnor (d125, d88, d90);
	buf (d126, d90);
	xnor (d127, d79, d86);
	xor (d128, d67, d89);
	not (d129, d18);
	xor (d130, d73, d86);
	and (d131, d74, d83);
	not (d132, d32);
	xor (d133, d70);
	xor (d134, d85, d91);
	nand (d135, d68, d69);
	nand (d136, d69, d88);
	not (d137, d79);
	nand (d138, d77, d88);
	xnor (d139, d71, d79);
	buf (d140, d46);
	buf (d141, d59);
	xor (d142, d71, d81);
	nand (d143, d77);
	or (d144, d69, d88);
	xnor (d145, d66, d80);
	or (d146, d71, d89);
	buf (d147, d13);
	xnor (d148, d83, d85);
	nand (d149, d84, d90);
	nor (d150, d83, d87);
	buf (d151, d56);
	or (d152, d67, d87);
	buf (d153, d7);
	xor (d154, d67, d71);
	nand (d155, d70, d90);
	and (d156, d84, d86);
	nand (d157, d70, d79);
	nand (d158, d69, d85);
	buf (d159, d21);
	nor (d160, d78, d83);
	xnor (d161, d127, d158);
	xor (d162, d133, d145);
	nand (d163, d114, d137);
	xor (d164, d97, d133);
	and (d165, d136, d153);
	xor (d166, d121, d160);
	and (d167, d121, d129);
	xor (d168, d104, d106);
	xnor (d169, d109, d135);
	and (d170, d121, d150);
	xor (d171, d94, d138);
	and (d172, d130, d158);
	nor (d173, d103, d143);
	nand (d174, d110, d121);
	not (d175, d62);
	xnor (d176, d110, d131);
	xnor (d177, d95, d139);
	xnor (d178, d101, d153);
	and (d179, d102, d114);
	buf (d180, d101);
	or (d181, d173, d174);
	or (d182, d175, d177);
	or (d183, d166, d177);
	not (d184, d146);
	buf (d185, d86);
	nand (d186, d171, d176);
	nand (d187, d161, d173);
	not (d188, d99);
	xnor (d189, d165, d173);
	and (d190, d165, d180);
	or (d191, d166, d180);
	nor (d192, d164, d171);
	and (d193, d172, d177);
	not (d194, d19);
	xnor (d195, d164, d167);
	not (d196, d56);
	xnor (d197, d166, d175);
	not (d198, d29);
	xor (d199, d164, d168);
	buf (d200, d49);
	nor (d201, d161, d172);
	buf (d202, d50);
	xnor (d203, d173, d179);
	or (d204, d173);
	nand (d205, d173, d177);
	nand (d206, d197);
	and (d207, d183, d202);
	xor (d208, d194, d196);
	xor (d209, d192, d197);
	or (d210, d198);
	or (d211, d182, d197);
	xnor (d212, d197, d202);
	buf (d213, d189);
	nor (d214, d183, d204);
	buf (d215, d142);
	nand (d216, d191, d199);
	and (d217, d181, d198);
	buf (d218, d199);
	buf (d219, d157);
	xor (d220, d190, d200);
	or (d221, d182, d194);
	nor (d222, d181, d203);
	buf (d223, d202);
	xnor (d224, d195);
	nor (d225, d182, d185);
	and (d226, d191, d200);
	and (d227, d192, d202);
	xnor (d228, d187, d196);
	and (d229, d187, d201);
	or (d230, d184, d194);
	xnor (d231, d192, d205);
	nand (d232, d192, d196);
	buf (d233, d191);
	nor (d234, d202, d203);
	nand (d235, d187, d201);
	xnor (d236, d185, d205);
	buf (d237, d4);
	or (d238, d202);
	or (d239, d190, d205);
	buf (d240, d198);
	nor (d241, d192, d201);
	nor (d242, d199, d200);
	xor (d243, d185, d188);
	not (d244, d22);
	nand (d245, d183, d201);
	buf (d246, d135);
	xnor (d247, d184, d205);
	not (d248, d164);
	nor (d249, d195, d203);
	xor (d250, d197, d205);
	xor (d251, d197, d203);
	buf (d252, d84);
	xor (d253, d191, d205);
	nor (d254, d186, d202);
	nor (d255, d187, d202);
	and (d256, d181, d183);
	nor (d257, d185, d197);
	xnor (d258, d197, d205);
	not (d259, d43);
	and (d260, d186, d205);
	nand (d261, d195, d200);
	not (d262, d172);
	xor (d263, d199, d201);
	xor (d264, d198);
	nand (d265, d190, d204);
	nor (d266, d195, d200);
	and (d267, d186, d187);
	nand (d268, d202, d205);
	nand (d269, d186, d195);
	or (d270, d186, d194);
	nor (d271, d187, d204);
	nand (d272, d192, d200);
	not (d273, d158);
	nor (d274, d189, d197);
	nor (d275, d196, d201);
	and (d276, d181, d192);
	nor (d277, d191, d204);
	xor (d278, d195, d199);
	xnor (d279, d184, d202);
	buf (d280, d82);
	buf (d281, d69);
	nor (d282, d189, d196);
	nand (d283, d182, d194);
	not (d284, d59);
	buf (d285, d205);
	buf (d286, d72);
	nor (d287, d199, d204);
	xnor (d288, d182, d188);
	and (d289, d185);
	xor (d290, d222, d243);
	nor (d291, d209, d262);
	xor (d292, d214, d235);
	not (d293, d176);
	nor (d294, d233, d278);
	xnor (d295, d231, d249);
	buf (d296, d61);
	nand (d297, d213, d277);
	xnor (d298, d233, d266);
	buf (d299, d238);
	not (d300, d141);
	xor (d301, d258, d270);
	or (d302, d207, d259);
	xor (d303, d251, d270);
	or (d304, d240, d246);
	nand (d305, d264, d278);
	and (d306, d215, d246);
	nor (d307, d227, d245);
	xor (d308, d215, d228);
	nor (d309, d250, d269);
	xor (d310, d218, d280);
	nand (d311, d233, d274);
	nor (d312, d213, d276);
	xor (d313, d213, d264);
	nand (d314, d212, d238);
	and (d315, d224, d284);
	nand (d316, d234, d273);
	not (d317, d42);
	xor (d318, d227, d274);
	xor (d319, d244, d262);
	nand (d320, d239, d265);
	xor (d321, d222, d237);
	nand (d322, d216, d223);
	not (d323, d25);
	buf (d324, d187);
	xor (d325, d274, d287);
	or (d326, d221, d229);
	or (d327, d247, d253);
	buf (d328, d171);
	and (d329, d224, d281);
	nand (d330, d237, d238);
	and (d331, d209, d223);
	nand (d332, d264, d278);
	buf (d333, d15);
	or (d334, d227, d266);
	nand (d335, d212, d239);
	nor (d336, d229, d235);
	or (d337, d238, d245);
	nand (d338, d231, d287);
	xor (d339, d209, d220);
	xnor (d340, d208, d225);
	nor (d341, d214, d244);
	buf (d342, d80);
	and (d343, d207, d216);
	not (d344, d264);
	or (d345, d254, d277);
	or (d346, d248, d249);
	and (d347, d230, d271);
	xor (d348, d245, d262);
	not (d349, d268);
	and (d350, d236, d287);
	or (d351, d208, d228);
	buf (d352, d57);
	not (d353, d337);
	or (d354, d314, d334);
	or (d355, d316, d336);
	xor (d356, d300, d335);
	buf (d357, d309);
	or (d358, d301, d316);
	and (d359, d291, d352);
	or (d360, d311, d352);
	or (d361, d310, d341);
	nor (d362, d307, d336);
	not (d363, d348);
	nor (d364, d327, d351);
	or (d365, d291, d319);
	xor (d366, d315, d317);
	xor (d367, d303, d308);
	or (d368, d293, d347);
	nor (d369, d291, d338);
	or (d370, d340, d348);
	buf (d371, d145);
	not (d372, d199);
	or (d373, d299, d334);
	and (d374, d350, d351);
	not (d375, d127);
	or (d376, d310, d314);
	and (d377, d312);
	nor (d378, d310, d325);
	nor (d379, d330, d342);
	buf (d380, d335);
	or (d381, d302, d329);
	nand (d382, d315, d334);
	or (d383, d324, d328);
	xor (d384, d339, d350);
	nor (d385, d299, d335);
	xor (d386, d341, d350);
	not (d387, d84);
	nand (d388, d292, d347);
	nor (d389, d323, d326);
	buf (d390, d138);
	xor (d391, d324, d333);
	or (d392, d301, d329);
	not (d393, d6);
	not (d394, d291);
	nand (d395, d322, d350);
	buf (d396, d228);
	nand (d397, d296, d340);
	not (d398, d125);
	buf (d399, d143);
	not (d400, d317);
	buf (d401, d47);
	nor (d402, d309, d319);
	and (d403, d334, d336);
	buf (d404, d55);
	nor (d405, d292, d305);
	nor (d406, d340, d341);
	nand (d407, d324, d334);
	xor (d408, d329, d340);
	not (d409, d220);
	or (d410, d325, d334);
	not (d411, d332);
	nand (d412, d320, d343);
	not (d413, d198);
	nand (d414, d350, d351);
	xor (d415, d322, d333);
	or (d416, d317, d352);
	xnor (d417, d300, d344);
	not (d418, d147);
	and (d419, d297, d336);
	buf (d420, d98);
	xnor (d421, d309, d316);
	xor (d422, d341);
	buf (d423, d239);
	xor (d424, d318, d335);
	nand (d425, d311, d350);
	or (d426, d299, d322);
	nor (d427, d290, d343);
	xor (d428, d323, d349);
	nor (d429, d291, d297);
	and (d430, d300, d301);
	xnor (d431, d296, d318);
	nand (d432, d306, d322);
	not (d433, d329);
	buf (d434, d129);
	xor (d435, d382, d413);
	and (d436, d361, d408);
	nand (d437, d366, d428);
	xor (d438, d377, d420);
	buf (d439, d333);
	xor (d440, d362, d428);
	not (d441, d189);
	xnor (d442, d356, d425);
	and (d443, d397, d433);
	or (d444, d387, d434);
	xnor (d445, d370, d402);
	xnor (d446, d364, d369);
	not (d447, d221);
	buf (d448, d314);
	xnor (d449, d375, d389);
	not (d450, d28);
	not (d451, d298);
	xor (d452, d372, d398);
	nor (d453, d369, d370);
	buf (d454, d58);
	nor (d455, d356, d415);
	xor (d456, d355, d411);
	buf (d457, d163);
	nor (d458, d357, d381);
	or (d459, d378, d398);
	xor (d460, d378, d427);
	and (d461, d359, d381);
	buf (d462, d78);
	xor (d463, d373, d424);
	and (d464, d363, d434);
	xor (d465, d419);
	nor (d466, d380, d388);
	xnor (d467, d371, d409);
	or (d468, d391, d404);
	or (d469, d391, d428);
	or (d470, d365, d412);
	and (d471, d383, d424);
	nand (d472, d385, d428);
	nand (d473, d354, d427);
	xor (d474, d379, d422);
	nand (d475, d364, d366);
	and (d476, d368, d418);
	nor (d477, d384, d393);
	buf (d478, d107);
	not (d479, d177);
	nor (d480, d390, d427);
	nor (d481, d360, d424);
	xor (d482, d386, d391);
	xnor (d483, d406, d427);
	not (d484, d45);
	nor (d485, d371);
	nor (d486, d361, d376);
	nor (d487, d368, d382);
	buf (d488, d71);
	xor (d489, d364, d421);
	and (d490, d390, d397);
	nor (d491, d358, d360);
	nor (d492, d383);
	buf (d493, d363);
	or (d494, d368, d386);
	and (d495, d363, d364);
	assign f1 = d485;
	assign f2 = d464;
	assign f3 = d462;
	assign f4 = d451;
	assign f5 = d438;
	assign f6 = d482;
	assign f7 = d482;
	assign f8 = d460;
	assign f9 = d440;
endmodule
