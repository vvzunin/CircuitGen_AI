module CCGRCG73( x0, x1, x2, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17, f18, f19 );

	input x0, x1, x2;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17, f18, f19;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309;

	and (d1, x0, x2);
	not (d2, x0);
	and (d3, x0);
	nand (d4, x0, x2);
	nor (d5, x1, x2);
	buf (d6, x2);
	not (d7, x1);
	buf (d8, x0);
	nand (d9, x0, x2);
	nor (d10, x0, x2);
	xor (d11, x1);
	xnor (d12, x0);
	not (d13, x2);
	nand (d14, x2);
	or (d15, x0, x1);
	xor (d16, x0, x1);
	xor (d17, x0, x1);
	xor (d18, x0, x2);
	nor (d19, x0, x2);
	xor (d20, x0);
	xnor (d21, x1, x2);
	and (d22, x1, x2);
	nand (d23, x0, x1);
	and (d24, x0, x1);
	and (d25, x1);
	and (d26, x1, x2);
	buf (d27, x1);
	xor (d28, x1, x2);
	or (d29, x1, x2);
	nor (d30, x0, x1);
	or (d31, x1);
	nand (d32, x1, x2);
	nand (d33, x0, x1);
	xnor (d34, x1);
	xor (d35, x0, x2);
	nor (d36, x2);
	nor (d37, x1, x2);
	or (d38, x0, x1);
	and (d39, x0, x1);
	xnor (d40, x2);
	xnor (d41, x0, x1);
	or (d42, x0);
	not (d43, d31);
	and (d44, d30, d42);
	nor (d45, d31, d41);
	and (d46, d19, d23);
	or (d47, d4, d31);
	not (d48, d33);
	buf (d49, d41);
	not (d50, d42);
	xor (d51, d2, d28);
	not (d52, d8);
	nand (d53, d15, d21);
	nand (d54, d14, d27);
	or (d55, d13, d38);
	not (d56, d22);
	xor (d57, d30, d36);
	xor (d58, d30, d39);
	nand (d59, d23, d29);
	nand (d60, d6, d15);
	xnor (d61, d7, d42);
	and (d62, d19, d36);
	buf (d63, d26);
	nand (d64, d16, d23);
	xnor (d65, d1, d41);
	buf (d66, d28);
	or (d67, d21, d42);
	nor (d68, d7, d27);
	nor (d69, d14, d20);
	or (d70, d5, d8);
	nand (d71, d2, d10);
	xnor (d72, d26, d38);
	xnor (d73, d6, d24);
	or (d74, d16, d29);
	nor (d75, d12, d25);
	nand (d76, d5, d39);
	buf (d77, d25);
	and (d78, d17, d21);
	xor (d79, d49, d72);
	nor (d80, d44, d67);
	or (d81, d46, d73);
	nor (d82, d49, d75);
	nor (d83, d54, d77);
	not (d84, d34);
	nand (d85, d58, d64);
	nand (d86, d61, d65);
	nand (d87, d58, d66);
	not (d88, d72);
	buf (d89, d48);
	nor (d90, d45, d55);
	nand (d91, d54, d70);
	and (d92, d47, d66);
	nor (d93, d71, d77);
	nand (d94, d57, d64);
	nand (d95, d43, d77);
	and (d96, d62, d75);
	and (d97, d61, d77);
	xnor (d98, d48, d69);
	buf (d99, d24);
	and (d100, d65, d68);
	nand (d101, d51, d54);
	and (d102, d50, d77);
	buf (d103, d59);
	not (d104, d20);
	xor (d105, d59, d60);
	nor (d106, d47, d48);
	and (d107, d76, d78);
	xor (d108, d49, d78);
	nand (d109, d58, d59);
	xor (d110, d50, d54);
	or (d111, d52, d72);
	or (d112, d49);
	nor (d113, d50, d53);
	or (d114, d57, d63);
	nor (d115, d50, d67);
	or (d116, d46, d74);
	not (d117, d13);
	buf (d118, d21);
	and (d119, d45, d49);
	xor (d120, d69, d71);
	or (d121, d66, d78);
	and (d122, d46, d64);
	and (d123, d46, d75);
	and (d124, d72, d76);
	and (d125, d44, d77);
	and (d126, d67, d77);
	and (d127, d49, d77);
	nand (d128, d48, d68);
	buf (d129, d51);
	and (d130, d56, d61);
	buf (d131, d15);
	nand (d132, d47, d65);
	and (d133, d62, d72);
	nor (d134, d58, d59);
	nand (d135, d69, d78);
	and (d136, d53, d66);
	not (d137, d62);
	xnor (d138, d46, d71);
	nor (d139, d70, d78);
	and (d140, d45, d69);
	nor (d141, d63, d76);
	xor (d142, d44);
	buf (d143, d22);
	or (d144, d46, d55);
	and (d145, d71, d78);
	buf (d146, d17);
	not (d147, d76);
	xor (d148, d69, d70);
	xor (d149, d47, d53);
	not (d150, d2);
	or (d151, d58, d72);
	xnor (d152, d54, d78);
	or (d153, d58, d69);
	nand (d154, d57, d76);
	or (d155, d49, d58);
	xnor (d156, d49, d57);
	nand (d157, d65, d68);
	and (d158, d44, d63);
	buf (d159, d7);
	xnor (d160, d60, d69);
	nand (d161, d62, d68);
	xor (d162, d50, d73);
	or (d163, d45, d57);
	nor (d164, d50, d63);
	xor (d165, d131, d138);
	nand (d166, d125, d138);
	buf (d167, d73);
	and (d168, d139, d142);
	nor (d169, d79, d108);
	nor (d170, d166, d169);
	not (d171, d102);
	nand (d172, d166);
	or (d173, d167);
	xor (d174, d166, d167);
	nand (d175, d167, d169);
	or (d176, d167, d168);
	not (d177, d97);
	not (d178, d111);
	nand (d179, d166, d167);
	xnor (d180, d165);
	or (d181, d166, d168);
	and (d182, d166, d168);
	and (d183, d165, d166);
	nor (d184, d168, d169);
	xor (d185, d167, d169);
	xor (d186, d165, d167);
	and (d187, d165, d167);
	nor (d188, d165, d168);
	xor (d189, d167, d169);
	xor (d190, d166, d169);
	nand (d191, d166, d168);
	or (d192, d165, d166);
	xor (d193, d165, d169);
	nor (d194, d165, d169);
	nor (d195, d166, d168);
	not (d196, d113);
	buf (d197, d164);
	not (d198, d112);
	not (d199, d57);
	xor (d200, d165, d166);
	nand (d201, d165, d168);
	not (d202, d74);
	buf (d203, d23);
	xor (d204, d165, d168);
	nand (d205, d167);
	and (d206, d165, d168);
	xnor (d207, d165, d169);
	xor (d208, d167);
	not (d209, d126);
	nand (d210, d168, d169);
	nor (d211, d165, d167);
	xor (d212, d166, d168);
	and (d213, d166, d169);
	not (d214, d18);
	or (d215, d166, d169);
	not (d216, d63);
	not (d217, d101);
	and (d218, d168, d169);
	not (d219, d82);
	xnor (d220, d165, d167);
	not (d221, d46);
	xnor (d222, d166, d168);
	xnor (d223, d167, d169);
	or (d224, d167, d169);
	nor (d225, d166, d167);
	buf (d226, d95);
	xor (d227, d167, d168);
	xnor (d228, d167, d168);
	or (d229, d168);
	and (d230, d167);
	and (d231, d166, d167);
	nand (d232, d166, d168);
	nand (d233, d173, d179);
	xor (d234, d203, d215);
	xor (d235, d192, d229);
	or (d236, d195, d219);
	or (d237, d187, d204);
	xnor (d238, d194, d218);
	nor (d239, d184, d200);
	nand (d240, d198, d227);
	xnor (d241, d209, d222);
	xnor (d242, d172, d222);
	nor (d243, d177, d189);
	xnor (d244, d193, d221);
	and (d245, d203, d220);
	nor (d246, d182, d194);
	or (d247, d171, d177);
	or (d248, d214, d231);
	xnor (d249, d174, d227);
	or (d250, d191);
	xnor (d251, d187, d212);
	and (d252, d218, d221);
	xnor (d253, d184, d229);
	xor (d254, d177, d185);
	buf (d255, d151);
	nand (d256, d188, d200);
	or (d257, d171, d193);
	not (d258, d88);
	and (d259, d185, d216);
	xor (d260, d196, d228);
	xor (d261, d176, d198);
	or (d262, d194, d219);
	buf (d263, d6);
	not (d264, d159);
	or (d265, d173, d197);
	xor (d266, d223, d231);
	xnor (d267, d190, d191);
	xnor (d268, d192, d205);
	and (d269, d176, d206);
	buf (d270, d42);
	xor (d271, d187, d189);
	xor (d272, d186, d211);
	xor (d273, d195, d207);
	nand (d274, d176, d224);
	not (d275, d145);
	xor (d276, d201, d203);
	nor (d277, d171, d178);
	xnor (d278, d171, d224);
	or (d279, d195, d220);
	or (d280, d201, d221);
	nand (d281, d176, d181);
	nor (d282, d205, d213);
	nand (d283, d187, d189);
	xnor (d284, d178, d204);
	not (d285, d136);
	or (d286, d199, d221);
	or (d287, d171, d198);
	not (d288, d24);
	xnor (d289, d174, d215);
	xnor (d290, d180, d232);
	nor (d291, d186, d194);
	and (d292, d209, d229);
	buf (d293, d35);
	xnor (d294, d186);
	nor (d295, d218, d229);
	xor (d296, d175, d189);
	xnor (d297, d224, d225);
	xor (d298, d171, d209);
	buf (d299, d19);
	xnor (d300, d173, d216);
	not (d301, d218);
	nand (d302, d200, d229);
	and (d303, d190, d203);
	nand (d304, d197, d224);
	nor (d305, d191, d221);
	xor (d306, d182, d217);
	nor (d307, d199, d215);
	or (d308, d181, d202);
	nand (d309, d202, d224);
	assign f1 = d248;
	assign f2 = d239;
	assign f3 = d250;
	assign f4 = d263;
	assign f5 = d289;
	assign f6 = d243;
	assign f7 = d239;
	assign f8 = d273;
	assign f9 = d255;
	assign f10 = d235;
	assign f11 = d293;
	assign f12 = d252;
	assign f13 = d280;
	assign f14 = d307;
	assign f15 = d241;
	assign f16 = d302;
	assign f17 = d270;
	assign f18 = d273;
	assign f19 = d254;
endmodule
