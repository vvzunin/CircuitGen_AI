// Benchmark "CCGRCG142" written by ABC on Tue Feb 13 20:52:06 2024

module CCGRCG142 ( 
    x0, x1, x2, x3, x4,
    f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16  );
  input  x0, x1, x2, x3, x4;
  output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15,
    f16;
  wire new_n22_, new_n23_, new_n24_, new_n25_, new_n26_, new_n27_, new_n28_,
    new_n29_, new_n30_, new_n31_, new_n33_, new_n34_, new_n35_, new_n36_,
    new_n37_, new_n38_, new_n39_, new_n40_, new_n41_, new_n43_, new_n44_,
    new_n45_, new_n47_, new_n48_, new_n49_, new_n50_, new_n51_, new_n52_,
    new_n53_, new_n55_, new_n59_, new_n60_, new_n61_, new_n62_, new_n63_,
    new_n65_, new_n66_, new_n67_, new_n70_, new_n71_, new_n72_, new_n75_,
    new_n76_, new_n77_, new_n78_, new_n79_;
  assign new_n22_ = x1 ^ x4;
  assign new_n23_ = ~x1;
  assign new_n24_ = ~new_n23_ | ~x2;
  assign new_n25_ = x2 | ~x1;
  assign new_n26_ = ~x0 | ~x3;
  assign new_n27_ = ~new_n26_;
  assign new_n28_ = ~x0;
  assign new_n29_ = ~x2;
  assign new_n30_ = ~x3;
  assign new_n31_ = ~new_n29_ | ~new_n28_ | (~x4 & ~new_n23_ & ~new_n30_);
  assign f1 = ~new_n27_ & ~new_n31_ & (~new_n22_ | ~new_n24_ | ~new_n25_);
  assign new_n33_ = ~x4;
  assign new_n34_ = ~x1 & ~new_n33_;
  assign new_n35_ = ~x4 | ~new_n29_ | ~x1;
  assign new_n36_ = ~x1 | ~x4;
  assign new_n37_ = ~new_n36_ | ~new_n24_ | ~new_n25_;
  assign new_n38_ = ~new_n37_ | ~new_n35_;
  assign new_n39_ = ~x0 & ~x2;
  assign new_n40_ = ~new_n28_ & ~new_n29_;
  assign new_n41_ = (~x1 & ~x3) | (~new_n39_ & ~new_n40_);
  assign f2 = ~new_n29_ & ~new_n34_ & ~new_n41_ & (~new_n38_ | ~new_n27_);
  assign new_n43_ = ~new_n39_;
  assign new_n44_ = ~new_n30_ | ~new_n33_;
  assign new_n45_ = ~new_n28_ | ~new_n23_;
  assign new_n47_ = ~x3 | ~x2 | ~new_n33_ | ~x1;
  assign new_n48_ = ~new_n43_ | (~new_n44_ & ~new_n47_);
  assign new_n49_ = ~new_n48_ | ~new_n27_;
  assign new_n50_ = ~new_n26_ | ~new_n43_ | (~new_n44_ & ~new_n47_);
  assign new_n51_ = new_n38_ & new_n50_ & new_n49_ & (new_n23_ | new_n30_);
  assign new_n52_ = ~x1 | ~x3;
  assign new_n53_ = (~new_n38_ | ~new_n52_) & (~new_n49_ | ~new_n50_);
  assign f3 = ~new_n53_ & ~new_n51_;
  assign new_n55_ = ~new_n29_ | (~new_n23_ & ~x4) | (~new_n26_ & ~new_n41_);
  assign f4 = ~new_n26_ | ~new_n33_ | ~new_n55_ | ~new_n29_;
  assign f5 = ~new_n43_ | ~new_n27_;
  assign f6 = ~new_n52_;
  assign new_n59_ = ~new_n28_ | ~x3;
  assign new_n60_ = ~new_n44_ | ~new_n59_;
  assign new_n61_ = ~new_n25_ | ~new_n33_;
  assign new_n62_ = ~new_n61_ | ~new_n24_;
  assign new_n63_ = new_n60_ ^ new_n62_;
  assign f9 = ~new_n31_ & ~new_n63_;
  assign new_n65_ = ~new_n36_ & (~new_n28_ | ~x2);
  assign new_n66_ = ~new_n33_ & ~new_n65_;
  assign new_n67_ = ~new_n23_ & ~x2 & (~new_n28_ | ~new_n30_ | ~new_n33_);
  assign f10 = ~new_n67_ | ~new_n66_;
  assign f11 = ~new_n31_ | (~x2 & ~new_n59_) | (~x3 & ~new_n48_);
  assign new_n70_ = ~new_n29_ | (~x4 & ~new_n23_) | (~new_n28_ & ~new_n30_);
  assign new_n71_ = ~new_n25_ | (~new_n29_ & ~new_n33_);
  assign new_n72_ = ~new_n70_ | ~new_n71_;
  assign f12 = ~new_n72_ & ~new_n39_ & ~new_n65_;
  assign new_n75_ = ~x0 & ~x2 & (~new_n30_ | ~new_n33_ | ~x1);
  assign new_n76_ = ~x2 | ~new_n28_ | ~new_n23_;
  assign new_n77_ = (new_n35_ & new_n37_) | (~new_n29_ & ~new_n45_);
  assign new_n78_ = ~new_n76_ | ~new_n77_ | ~new_n75_;
  assign new_n79_ = ~new_n78_ | ~new_n31_;
  assign f14 = ~new_n79_ | (~new_n55_ & ~new_n78_);
  assign f15 = ~new_n71_ & (~new_n33_ | ~new_n52_);
  assign f16 = ~new_n39_ | ~new_n30_;
  assign f13 = 1'b1;
  assign f7 = ~new_n53_ & ~new_n51_;
  assign f8 = ~new_n52_;
endmodule


