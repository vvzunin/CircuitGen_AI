module CCGRCG78( x0, x1, x2, x3, f1, f2, f3 );

	input x0, x1, x2, x3;
	output f1, f2, f3;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314, d315, d316, d317, d318, d319, d320, d321, d322, d323, d324, d325, d326, d327, d328, d329, d330, d331, d332, d333, d334, d335, d336, d337, d338, d339, d340, d341, d342, d343, d344, d345, d346, d347, d348, d349, d350, d351, d352, d353, d354, d355, d356, d357, d358, d359, d360, d361, d362, d363, d364, d365, d366, d367, d368, d369, d370, d371, d372, d373, d374, d375, d376, d377, d378, d379, d380, d381, d382, d383, d384, d385, d386, d387, d388, d389, d390, d391, d392, d393, d394, d395, d396, d397, d398, d399, d400, d401, d402, d403, d404, d405, d406;

	buf (d1, x1);
	nor (d2, x0, x2);
	and (d3, x2, x3);
	or (d4, x1);
	nand (d5, x0, x1);
	xnor (d6, x1, x2);
	nor (d7, x1, x2);
	xnor (d8, x3);
	not (d9, x0);
	and (d10, x0, x3);
	nand (d11, x0, x3);
	or (d12, x1, x2);
	nor (d13, x1);
	xnor (d14, x1, x3);
	and (d15, x1, x2);
	and (d16, x1, x2);
	xor (d17, x0, x1);
	nor (d18, x1, x3);
	xnor (d19, x2);
	nand (d20, x1, x3);
	xnor (d21, x0, x3);
	xnor (d22, x0, x1);
	xnor (d23, x1, x2);
	not (d24, x1);
	buf (d25, x3);
	and (d26, x0, x2);
	xor (d27, x2);
	nand (d28, x0);
	nor (d29, x0, x2);
	nor (d30, x3);
	buf (d31, x2);
	nor (d32, x0, x1);
	xnor (d33, x2, x3);
	xor (d34, x1, x2);
	xor (d35, x2, x3);
	not (d36, x3);
	nand (d37, x2, x3);
	xor (d38, x0, x2);
	or (d39, x0, x2);
	xor (d40, x0, x3);
	or (d41, x1, x3);
	nand (d42, x2);
	xor (d43, x0);
	nand (d44, x1, x2);
	nor (d45, x1, x2);
	and (d46, x0, x2);
	nand (d47, x0, x2);
	nor (d48, d5, d20);
	xor (d49, d36, d45);
	or (d50, d2, d13);
	buf (d51, x0);
	xor (d52, d24, d26);
	buf (d53, d27);
	xor (d54, d4, d26);
	xor (d55, d19, d29);
	and (d56, d22, d30);
	nand (d57, d3, d7);
	xor (d58, d16, d46);
	nor (d59, d11, d38);
	xor (d60, d27, d29);
	not (d61, d38);
	nor (d62, d14, d36);
	xnor (d63, d21, d46);
	xnor (d64, d6, d44);
	not (d65, d31);
	nand (d66, d3, d11);
	and (d67, d22, d23);
	not (d68, d7);
	or (d69, d40, d41);
	buf (d70, d20);
	buf (d71, d33);
	or (d72, d19, d34);
	buf (d73, d1);
	or (d74, d18, d20);
	or (d75, d19, d25);
	nand (d76, d3, d21);
	nor (d77, d26, d32);
	buf (d78, d17);
	not (d79, d17);
	xor (d80, d7, d42);
	or (d81, d8, d42);
	or (d82, d30, d31);
	xnor (d83, d3, d30);
	buf (d84, d37);
	xnor (d85, d2, d34);
	or (d86, d15, d17);
	xor (d87, d29, d33);
	nand (d88, d18, d43);
	xnor (d89, d8, d22);
	nor (d90, d25, d47);
	nand (d91, d7, d11);
	or (d92, d39, d47);
	not (d93, d6);
	xnor (d94, d10, d26);
	nand (d95, d2, d36);
	buf (d96, d45);
	nand (d97, d22, d40);
	xor (d98, d26, d41);
	or (d99, d10, d15);
	or (d100, d34);
	nor (d101, d26, d33);
	and (d102, d11, d25);
	nor (d103, d29, d44);
	nor (d104, d1, d42);
	xnor (d105, d17, d26);
	xor (d106, d1, d24);
	nand (d107, d10, d34);
	or (d108, d7, d34);
	buf (d109, d18);
	and (d110, d72, d78);
	nand (d111, d70, d96);
	not (d112, d19);
	xor (d113, d107, d108);
	not (d114, d101);
	nor (d115, d51, d105);
	and (d116, d54, d103);
	not (d117, d60);
	not (d118, d55);
	or (d119, d91, d97);
	buf (d120, d91);
	and (d121, d57, d68);
	xor (d122, d68, d79);
	not (d123, d105);
	nand (d124, d50, d52);
	nor (d125, d61, d78);
	or (d126, d49, d74);
	xnor (d127, d65, d72);
	buf (d128, d26);
	or (d129, d60, d94);
	nand (d130, d67, d72);
	nand (d131, d82, d106);
	buf (d132, d53);
	not (d133, d44);
	or (d134, d77, d109);
	nand (d135, d122, d130);
	nand (d136, d124, d130);
	and (d137, d112, d122);
	nor (d138, d112, d119);
	and (d139, d114, d123);
	not (d140, d107);
	and (d141, d111, d130);
	or (d142, d115, d133);
	xor (d143, d110, d134);
	or (d144, d120, d121);
	and (d145, d123, d130);
	xor (d146, d125, d133);
	xor (d147, d114, d124);
	nand (d148, d117, d131);
	or (d149, d110, d118);
	nor (d150, d118, d121);
	nor (d151, d126);
	nand (d152, d117, d118);
	xor (d153, d118, d124);
	xnor (d154, d114, d129);
	xnor (d155, d121, d134);
	nand (d156, d116, d131);
	xor (d157, d115, d126);
	and (d158, d114, d126);
	nand (d159, d130, d134);
	or (d160, d130, d134);
	xnor (d161, d127, d128);
	or (d162, d110, d125);
	nor (d163, d112, d119);
	or (d164, d110, d130);
	nand (d165, d116, d127);
	or (d166, d110, d117);
	or (d167, d114, d126);
	nor (d168, d112, d131);
	buf (d169, d49);
	nor (d170, d113, d133);
	or (d171, d120, d127);
	xor (d172, d111, d117);
	nand (d173, d129, d134);
	or (d174, d110, d129);
	nand (d175, d110, d122);
	xnor (d176, d118, d125);
	xor (d177, d123, d125);
	xnor (d178, d111, d122);
	not (d179, d37);
	nor (d180, d111, d124);
	nor (d181, d125, d129);
	and (d182, d111, d122);
	xnor (d183, d122, d128);
	nor (d184, d110, d130);
	not (d185, d22);
	buf (d186, d50);
	xor (d187, d113, d121);
	buf (d188, d56);
	nand (d189, d120, d127);
	nand (d190, d116, d133);
	and (d191, d120, d122);
	buf (d192, d51);
	not (d193, d51);
	buf (d194, d68);
	buf (d195, d21);
	nor (d196, d111, d130);
	or (d197, d124);
	nor (d198, d124, d130);
	nor (d199, d111, d112);
	xnor (d200, d110, d127);
	xnor (d201, d125, d129);
	nor (d202, d117, d128);
	nor (d203, d124, d125);
	buf (d204, d124);
	buf (d205, d133);
	buf (d206, d65);
	nand (d207, d113, d132);
	nand (d208, d117, d125);
	nand (d209, d157, d191);
	not (d210, d35);
	nand (d211, d140, d167);
	and (d212, d182, d193);
	nand (d213, d159, d174);
	nor (d214, d156, d198);
	nor (d215, d163, d195);
	nor (d216, d158, d177);
	nor (d217, d151, d198);
	and (d218, d135, d177);
	or (d219, d165, d180);
	xnor (d220, d149, d184);
	not (d221, d40);
	buf (d222, d5);
	nand (d223, d138, d173);
	xnor (d224, d155, d184);
	nor (d225, d143, d207);
	xor (d226, d170, d188);
	xor (d227, d158, d175);
	xor (d228, d152, d170);
	and (d229, d146, d155);
	not (d230, d103);
	and (d231, d142, d195);
	nand (d232, d156, d177);
	and (d233, d135, d194);
	buf (d234, d96);
	and (d235, d140, d207);
	or (d236, d135, d199);
	nand (d237, d150, d193);
	nor (d238, d194, d198);
	buf (d239, d177);
	xor (d240, d177, d205);
	nor (d241, d141, d160);
	and (d242, d154, d192);
	nor (d243, d158, d167);
	not (d244, d207);
	or (d245, d194, d205);
	xor (d246, d186, d188);
	nor (d247, d139, d153);
	xnor (d248, d138, d197);
	nand (d249, d152, d157);
	and (d250, d199, d207);
	not (d251, d9);
	buf (d252, d38);
	nand (d253, d189, d195);
	xor (d254, d135, d163);
	or (d255, d153, d207);
	and (d256, d170, d204);
	xnor (d257, d147, d207);
	and (d258, d150, d188);
	or (d259, d148, d202);
	xor (d260, d175, d184);
	and (d261, d165, d170);
	not (d262, d197);
	or (d263, d147, d182);
	or (d264, d172, d193);
	and (d265, d148, d155);
	not (d266, d33);
	and (d267, d140, d161);
	buf (d268, d40);
	or (d269, d219, d235);
	nand (d270, d226, d254);
	nor (d271, d227, d228);
	nand (d272, d258, d265);
	xnor (d273, d222, d230);
	xor (d274, d209, d223);
	xor (d275, d240, d258);
	and (d276, d258, d266);
	xnor (d277, d234, d236);
	and (d278, d234, d237);
	xor (d279, d226, d254);
	not (d280, d100);
	buf (d281, d235);
	xor (d282, d220, d233);
	xor (d283, d225, d234);
	buf (d284, d237);
	nor (d285, d215, d239);
	not (d286, d132);
	or (d287, d237, d262);
	buf (d288, d113);
	xor (d289, d220, d240);
	not (d290, d64);
	or (d291, d211, d251);
	nand (d292, d247, d255);
	nand (d293, d250, d263);
	nand (d294, d214, d243);
	buf (d295, d69);
	or (d296, d216, d248);
	nor (d297, d209, d246);
	xor (d298, d227, d240);
	nor (d299, d253, d258);
	buf (d300, d111);
	or (d301, d245, d258);
	and (d302, d226, d252);
	or (d303, d211, d266);
	nor (d304, d218, d249);
	xor (d305, d219, d255);
	and (d306, d216, d239);
	nor (d307, d225, d246);
	xor (d308, d239, d266);
	or (d309, d244, d265);
	xnor (d310, d215, d260);
	or (d311, d210, d214);
	or (d312, d213, d255);
	nand (d313, d219, d247);
	not (d314, d267);
	xnor (d315, d209, d218);
	xnor (d316, d234, d235);
	or (d317, d213, d243);
	buf (d318, d83);
	or (d319, d223, d253);
	or (d320, d254, d267);
	xor (d321, d248, d266);
	buf (d322, d120);
	xor (d323, d226, d258);
	xor (d324, d217, d263);
	xor (d325, d250, d261);
	xor (d326, d234, d240);
	and (d327, d249, d259);
	not (d328, d245);
	or (d329, d223, d237);
	not (d330, d85);
	and (d331, d211, d239);
	or (d332, d216, d218);
	not (d333, d141);
	nand (d334, d252, d262);
	buf (d335, d29);
	and (d336, d290, d295);
	buf (d337, d247);
	nand (d338, d274, d293);
	or (d339, d311, d330);
	buf (d340, d230);
	nor (d341, d314, d334);
	and (d342, d279, d329);
	xnor (d343, d271, d295);
	buf (d344, d52);
	xor (d345, d290, d327);
	or (d346, d292, d314);
	not (d347, d262);
	nand (d348, d302, d316);
	or (d349, d280, d299);
	nor (d350, d278, d301);
	buf (d351, d323);
	or (d352, d292, d297);
	not (d353, d29);
	and (d354, d295, d327);
	xor (d355, d311, d312);
	not (d356, d227);
	not (d357, d66);
	not (d358, d34);
	and (d359, d277, d295);
	xnor (d360, d302, d326);
	xor (d361, d286, d329);
	nand (d362, d292, d314);
	nor (d363, d319, d325);
	xnor (d364, d282, d316);
	buf (d365, d312);
	nand (d366, d322);
	nor (d367, d282, d318);
	buf (d368, d207);
	buf (d369, d99);
	nand (d370, d308, d313);
	xor (d371, d343, d363);
	or (d372, d348, d368);
	nor (d373, d350, d355);
	buf (d374, d366);
	nand (d375, d342, d356);
	buf (d376, d314);
	xor (d377, d359, d360);
	and (d378, d344, d360);
	xnor (d379, d353, d367);
	nor (d380, d339, d343);
	xnor (d381, d346, d364);
	not (d382, d58);
	buf (d383, d179);
	xnor (d384, d337, d357);
	nand (d385, d346, d359);
	xor (d386, d347, d352);
	and (d387, d353, d370);
	nor (d388, d353, d368);
	xnor (d389, d336, d352);
	nand (d390, d340, d360);
	xor (d391, d345, d357);
	buf (d392, d59);
	or (d393, d335, d366);
	xnor (d394, d341, d364);
	buf (d395, d154);
	nand (d396, d342, d368);
	xor (d397, d346, d350);
	nand (d398, d346, d351);
	nand (d399, d342, d370);
	nor (d400, d367, d368);
	or (d401, d340, d346);
	xor (d402, d347, d362);
	nand (d403, d358, d368);
	xor (d404, d339, d350);
	xnor (d405, d362, d363);
	not (d406, d82);
	assign f1 = d401;
	assign f2 = d372;
	assign f3 = d387;
endmodule
