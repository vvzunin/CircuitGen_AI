module CCGRCG39( x0, x1, x2, x3, x4, x5, x6, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12 );

	input x0, x1, x2, x3, x4, x5, x6;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314, d315, d316, d317, d318, d319, d320, d321, d322, d323, d324, d325, d326, d327, d328, d329, d330, d331, d332, d333, d334, d335, d336, d337, d338, d339, d340, d341, d342, d343, d344, d345, d346, d347, d348, d349, d350, d351, d352, d353, d354, d355, d356, d357, d358, d359, d360, d361, d362, d363, d364, d365, d366, d367, d368, d369, d370, d371, d372, d373, d374, d375, d376, d377, d378, d379, d380, d381, d382, d383, d384, d385, d386, d387, d388, d389, d390, d391, d392, d393, d394, d395, d396, d397, d398, d399, d400, d401, d402, d403, d404, d405, d406, d407, d408, d409, d410, d411, d412, d413, d414, d415, d416, d417, d418, d419, d420, d421, d422, d423, d424, d425, d426, d427, d428, d429, d430, d431, d432, d433, d434, d435, d436, d437, d438, d439, d440, d441, d442, d443, d444, d445, d446, d447, d448, d449, d450, d451, d452, d453, d454, d455, d456, d457, d458, d459, d460, d461, d462, d463, d464, d465, d466, d467, d468, d469, d470, d471, d472, d473, d474, d475, d476, d477, d478, d479, d480, d481, d482, d483, d484, d485, d486, d487, d488, d489, d490, d491, d492, d493, d494, d495, d496, d497, d498, d499, d500, d501, d502, d503, d504, d505, d506, d507, d508, d509, d510, d511, d512, d513, d514, d515, d516, d517, d518, d519, d520, d521, d522, d523, d524, d525, d526, d527, d528, d529, d530, d531, d532, d533, d534, d535, d536, d537, d538, d539, d540, d541, d542, d543, d544, d545, d546, d547, d548, d549, d550, d551, d552, d553, d554, d555, d556, d557, d558, d559, d560, d561, d562, d563, d564, d565, d566, d567, d568, d569, d570, d571, d572, d573, d574, d575, d576, d577, d578, d579, d580, d581, d582, d583, d584, d585, d586, d587, d588, d589, d590, d591, d592, d593, d594, d595, d596, d597, d598, d599, d600, d601, d602, d603, d604, d605, d606, d607, d608, d609, d610, d611, d612, d613, d614, d615, d616, d617, d618, d619, d620, d621, d622, d623, d624, d625, d626, d627, d628, d629, d630, d631, d632, d633, d634, d635, d636, d637, d638, d639, d640, d641, d642, d643, d644, d645, d646, d647, d648, d649, d650, d651, d652, d653, d654, d655, d656, d657, d658, d659, d660, d661, d662, d663, d664, d665, d666, d667, d668, d669, d670, d671, d672, d673, d674, d675, d676, d677, d678, d679, d680, d681, d682, d683, d684, d685, d686, d687, d688, d689, d690, d691, d692, d693, d694, d695, d696, d697, d698, d699, d700, d701, d702, d703, d704, d705, d706, d707, d708, d709, d710, d711, d712, d713, d714, d715, d716, d717, d718, d719, d720, d721, d722, d723, d724, d725, d726, d727, d728, d729, d730, d731, d732, d733, d734, d735, d736, d737, d738, d739, d740, d741, d742, d743, d744, d745, d746, d747, d748, d749, d750, d751, d752, d753, d754, d755, d756, d757, d758, d759, d760, d761, d762, d763, d764, d765, d766, d767, d768, d769, d770, d771, d772, d773, d774, d775, d776, d777, d778, d779, d780, d781, d782, d783, d784, d785, d786, d787, d788, d789, d790, d791, d792, d793, d794, d795, d796, d797, d798, d799, d800, d801, d802, d803, d804, d805, d806, d807, d808, d809, d810, d811, d812, d813, d814, d815, d816, d817, d818, d819, d820, d821, d822, d823, d824, d825, d826, d827, d828, d829, d830, d831, d832, d833, d834, d835;

	nand ( d1, x2, x3);
	buf ( d2, x5);
	nand ( d3, x5);
	nor ( d4, x0, x1);
	or ( d5, x1, x3);
	xnor ( d6, x3, x6);
	nor ( d7, x1, x4);
	and ( d8, x1, x2);
	xor ( d9, x3, x5);
	and ( d10, x0, x2);
	and ( d11, x0, x1);
	nand ( d12, x5, x6);
	not ( d13, x0);
	nand ( d14, x2, x6);
	xor ( d15, x4, x6);
	nor ( d16, x1, x4);
	xnor ( d17, x2, x3);
	nor ( d18, x0, x5);
	or ( d19, x0, x3);
	not ( d20, x4);
	buf ( d21, x0);
	or ( d22, x0, x4);
	nand ( d23, x0, x6);
	nor ( d24, x0, x1);
	not ( d25, x2);
	or ( d26, x2);
	xnor ( d27, x5);
	buf ( d28, x6);
	not ( d29, x5);
	xor ( d30, x3, x6);
	or ( d31, x2, x4);
	and ( d32, x2, x4);
	xor ( d33, x1, x5);
	nand ( d34, x3);
	not ( d35, x6);
	xnor ( d36, x0, x3);
	and ( d37, x4, x6);
	or ( d38, x3, x5);
	buf ( d39, x2);
	xor ( d40, x0);
	and ( d41, d32, d39);
	not ( d42, d9);
	not ( d43, x1);
	and ( d44, d7, d38);
	buf ( d45, d20);
	buf ( d46, d4);
	not ( d47, d36);
	or ( d48, d41, d43);
	xnor ( d49, d45, d46);
	buf ( d50, d24);
	not ( d51, d26);
	xnor ( d52, d42, d46);
	buf ( d53, d44);
	and ( d54, d45, d46);
	or ( d55, d42, d46);
	buf ( d56, d19);
	nor ( d57, d42, d46);
	xnor ( d58, d42, d45);
	buf ( d59, d3);
	buf ( d60, x3);
	or ( d61, d43, d46);
	nor ( d62, d42, d46);
	or ( d63, d44, d45);
	xor ( d64, d42, d44);
	nor ( d65, d41, d45);
	buf ( d66, d29);
	and ( d67, d44, d46);
	and ( d68, d41, d43);
	xnor ( d69, d41, d42);
	buf ( d70, d7);
	not ( d71, d3);
	and ( d72, d41, d42);
	and ( d73, d45, d46);
	and ( d74, d42, d44);
	nor ( d75, d45, d46);
	nor ( d76, d41, d44);
	and ( d77, d41, d45);
	buf ( d78, d12);
	and ( d79, d44);
	xor ( d80, d44, d46);
	not ( d81, d1);
	nor ( d82, d43, d46);
	nand ( d83, d41, d45);
	xor ( d84, d41, d45);
	or ( d85, d41, d44);
	not ( d86, d5);
	or ( d87, d41, d44);
	xnor ( d88, d43, d44);
	or ( d89, d51, d58);
	nand ( d90, d55);
	not ( d91, d16);
	xor ( d92, d55, d79);
	xnor ( d93, d49, d78);
	not ( d94, d33);
	xnor ( d95, d78, d84);
	or ( d96, d62, d73);
	xor ( d97, d58, d76);
	or ( d98, d60, d64);
	nand ( d99, d74, d75);
	not ( d100, d23);
	buf ( d101, d34);
	buf ( d102, d86);
	and ( d103, d62, d74);
	xnor ( d104, d64, d87);
	xnor ( d105, d55, d80);
	buf ( d106, d71);
	nand ( d107, d61, d73);
	nor ( d108, d68, d82);
	nor ( d109, d59, d65);
	xor ( d110, d51, d78);
	buf ( d111, d74);
	and ( d112, d51, d62);
	nand ( d113, d82);
	and ( d114, d109, d111);
	and ( d115, d96, d113);
	or ( d116, d89, d109);
	nand ( d117, d93, d104);
	and ( d118, d89, d95);
	nand ( d119, d95, d108);
	or ( d120, d105, d113);
	xor ( d121, d97, d113);
	not ( d122, d15);
	nor ( d123, d100, d113);
	or ( d124, d100, d106);
	xor ( d125, d99, d107);
	and ( d126, d91, d100);
	and ( d127, d106, d112);
	or ( d128, d97, d104);
	nand ( d129, d91, d95);
	not ( d130, d22);
	xnor ( d131, d110, d113);
	xor ( d132, d105, d113);
	nor ( d133, d94, d105);
	xnor ( d134, d96, d110);
	buf ( d135, d83);
	xor ( d136, d95, d107);
	not ( d137, d21);
	xnor ( d138, d97, d106);
	xnor ( d139, d93, d107);
	nor ( d140, d104, d108);
	xor ( d141, d97, d112);
	xnor ( d142, d96, d112);
	nor ( d143, d115, d141);
	nor ( d144, d114, d132);
	nor ( d145, d132, d137);
	buf ( d146, d111);
	nor ( d147, d126, d139);
	not ( d148, d103);
	or ( d149, d132, d136);
	not ( d150, d142);
	buf ( d151, d11);
	nand ( d152, d114, d136);
	xnor ( d153, d127, d130);
	xnor ( d154, d120, d141);
	nor ( d155, d118, d123);
	nand ( d156, d115, d127);
	or ( d157, d122, d129);
	and ( d158, d119, d122);
	nand ( d159, d126, d138);
	nand ( d160, d116, d126);
	xor ( d161, d115, d116);
	xor ( d162, d137, d139);
	not ( d163, d141);
	nor ( d164, d123, d142);
	buf ( d165, d46);
	not ( d166, d109);
	and ( d167, d119, d136);
	nor ( d168, d114, d119);
	and ( d169, d116, d119);
	not ( d170, d139);
	and ( d171, d138, d140);
	and ( d172, d130, d131);
	nor ( d173, d114, d115);
	nand ( d174, d126, d140);
	and ( d175, d126, d137);
	xor ( d176, d127, d134);
	xnor ( d177, d116, d128);
	and ( d178, d117, d136);
	xnor ( d179, d126, d134);
	xor ( d180, d137, d140);
	buf ( d181, d141);
	xor ( d182, d117, d124);
	nor ( d183, d130);
	nor ( d184, d114, d118);
	nand ( d185, d124, d129);
	and ( d186, d114, d137);
	xnor ( d187, d115, d142);
	not ( d188, d44);
	xnor ( d189, d117, d131);
	nand ( d190, d124, d137);
	or ( d191, d150, d151);
	buf ( d192, d156);
	nand ( d193, d154, d164);
	xnor ( d194, d147, d149);
	xor ( d195, d150, d160);
	xnor ( d196, d153, d164);
	or ( d197, d169, d171);
	xnor ( d198, d148, d166);
	buf ( d199, d164);
	nand ( d200, d155, d156);
	nand ( d201, d167, d176);
	xnor ( d202, d155, d158);
	xnor ( d203, d184, d189);
	or ( d204, d160, d162);
	and ( d205, d150, d155);
	nor ( d206, d170, d171);
	nor ( d207, d154, d167);
	or ( d208, d149, d164);
	buf ( d209, d75);
	nand ( d210, d157, d169);
	nand ( d211, d193, d197);
	or ( d212, d191, d203);
	nor ( d213, d204, d207);
	nor ( d214, d191, d194);
	not ( d215, x3);
	and ( d216, d200, d204);
	buf ( d217, d198);
	buf ( d218, d200);
	xnor ( d219, d206);
	xnor ( d220, d196, d198);
	nor ( d221, d191, d201);
	not ( d222, d47);
	and ( d223, d202, d208);
	xnor ( d224, d202, d210);
	buf ( d225, x1);
	not ( d226, d145);
	or ( d227, d214, d216);
	not ( d228, d169);
	xor ( d229, d215, d221);
	nand ( d230, d217, d219);
	nor ( d231, d218, d225);
	not ( d232, d160);
	not ( d233, d154);
	and ( d234, d212, d225);
	nand ( d235, d220, d224);
	buf ( d236, d196);
	buf ( d237, d185);
	xnor ( d238, d212, d223);
	nand ( d239, d212, d223);
	xor ( d240, d216, d219);
	not ( d241, d89);
	nand ( d242, d212, d218);
	nand ( d243, d213, d220);
	nand ( d244, d219, d221);
	or ( d245, d214, d223);
	xnor ( d246, d214, d223);
	and ( d247, d213, d220);
	and ( d248, d213, d223);
	xor ( d249, d212, d219);
	not ( d250, d113);
	and ( d251, d236, d248);
	and ( d252, d237, d250);
	or ( d253, d244, d248);
	nor ( d254, d251, d253);
	xnor ( d255, d252);
	xor ( d256, d252, d253);
	xor ( d257, d251);
	or ( d258, d253);
	nand ( d259, d251, d253);
	xnor ( d260, d251, d253);
	xor ( d261, d252, d253);
	and ( d262, d251);
	not ( d263, d218);
	nor ( d264, d251);
	not ( d265, d84);
	xor ( d266, d251, d253);
	and ( d267, d252, d253);
	nor ( d268, d252);
	nand ( d269, d251, d253);
	nor ( d270, d251, d252);
	and ( d271, d251, d252);
	or ( d272, d251, d253);
	nor ( d273, d252, d253);
	or ( d274, d251);
	nand ( d275, d253);
	buf ( d276, d239);
	and ( d277, d253);
	xnor ( d278, d251, d253);
	not ( d279, d90);
	not ( d280, d194);
	and ( d281, d252, d253);
	xnor ( d282, d252, d253);
	buf ( d283, d272);
	not ( d284, d120);
	nor ( d285, d257, d280);
	xnor ( d286, d262, d271);
	or ( d287, d255, d275);
	nand ( d288, d258, d274);
	xnor ( d289, d254, d259);
	xor ( d290, d264, d280);
	buf ( d291, d77);
	or ( d292, d254, d255);
	nand ( d293, d255, d258);
	nand ( d294, d262, d274);
	buf ( d295, d23);
	xor ( d296, d257, d277);
	not ( d297, d210);
	and ( d298, d254, d276);
	and ( d299, d255, d268);
	nor ( d300, d256, d257);
	xnor ( d301, d260, d261);
	nand ( d302, d262, d267);
	nor ( d303, d267, d273);
	and ( d304, d264, d281);
	xor ( d305, d269, d282);
	or ( d306, d267, d281);
	xnor ( d307, d267, d277);
	nor ( d308, d270, d279);
	nor ( d309, d268, d270);
	nand ( d310, d258, d261);
	xor ( d311, d273, d278);
	nor ( d312, d274, d281);
	or ( d313, d258, d271);
	and ( d314, d258, d266);
	xor ( d315, d268, d276);
	and ( d316, d269, d276);
	buf ( d317, d186);
	nor ( d318, d268, d270);
	or ( d319, d258, d264);
	or ( d320, d274, d275);
	nor ( d321, d284, d320);
	nand ( d322, d289, d315);
	xnor ( d323, d310, d320);
	xnor ( d324, d307, d308);
	or ( d325, d296, d301);
	xor ( d326, d286, d318);
	buf ( d327, d52);
	xnor ( d328, d285, d316);
	nand ( d329, d288, d299);
	nor ( d330, d285, d305);
	xor ( d331, d301, d317);
	xnor ( d332, d298, d299);
	buf ( d333, d163);
	xor ( d334, d288, d319);
	nand ( d335, d305, d308);
	nor ( d336, d305, d308);
	and ( d337, d283, d284);
	nor ( d338, d302, d312);
	xnor ( d339, d285, d298);
	not ( d340, d147);
	buf ( d341, d150);
	nand ( d342, d311, d318);
	nor ( d343, d292, d293);
	nor ( d344, d310, d311);
	xor ( d345, d296, d303);
	nor ( d346, d290, d301);
	not ( d347, d54);
	buf ( d348, d16);
	xnor ( d349, d302, d317);
	nand ( d350, d287, d301);
	xor ( d351, d294, d312);
	nand ( d352, d294, d315);
	xor ( d353, d284, d300);
	buf ( d354, d67);
	not ( d355, d167);
	or ( d356, d285, d293);
	buf ( d357, d292);
	or ( d358, d283, d308);
	and ( d359, d294, d317);
	and ( d360, d305, d320);
	xor ( d361, d286, d309);
	nor ( d362, d283, d289);
	nor ( d363, d292, d312);
	and ( d364, d295, d307);
	xor ( d365, d287, d305);
	xnor ( d366, d291, d315);
	buf ( d367, d72);
	nor ( d368, d294, d307);
	buf ( d369, d136);
	and ( d370, d331, d351);
	nor ( d371, d321, d368);
	xor ( d372, d352, d364);
	buf ( d373, d273);
	or ( d374, d335, d349);
	not ( d375, d318);
	xor ( d376, d332, d365);
	xnor ( d377, d324, d363);
	nor ( d378, d339, d364);
	xor ( d379, d357, d363);
	not ( d380, d12);
	xor ( d381, d352, d362);
	or ( d382, d332, d347);
	and ( d383, d337, d350);
	nor ( d384, d338, d341);
	nand ( d385, d323, d363);
	nor ( d386, d329, d354);
	buf ( d387, d15);
	nor ( d388, d347, d351);
	not ( d389, d315);
	nor ( d390, d328, d368);
	buf ( d391, d2);
	nor ( d392, d323, d336);
	and ( d393, d333, d349);
	xnor ( d394, d343, d345);
	and ( d395, d327, d336);
	nor ( d396, d336, d341);
	xor ( d397, d350, d362);
	buf ( d398, d132);
	nand ( d399, d360, d368);
	not ( d400, d243);
	not ( d401, d197);
	not ( d402, d339);
	nor ( d403, d322, d365);
	xor ( d404, d322, d343);
	xor ( d405, d325, d353);
	buf ( d406, d187);
	not ( d407, d337);
	buf ( d408, d364);
	nor ( d409, d347, d353);
	or ( d410, d392, d399);
	xor ( d411, d377, d399);
	nand ( d412, d372, d393);
	nor ( d413, d375);
	not ( d414, d88);
	nor ( d415, d374, d384);
	and ( d416, d384, d397);
	xor ( d417, d374, d401);
	xor ( d418, d369, d381);
	xor ( d419, d380, d389);
	buf ( d420, d129);
	and ( d421, d372, d377);
	buf ( d422, d276);
	or ( d423, d380, d389);
	xor ( d424, d374, d378);
	xor ( d425, d378);
	buf ( d426, d144);
	and ( d427, d394, d402);
	buf ( d428, d275);
	or ( d429, d382, d405);
	buf ( d430, d303);
	nor ( d431, d414, d415);
	and ( d432, d419);
	buf ( d433, d84);
	xnor ( d434, d424, d427);
	buf ( d435, d226);
	nor ( d436, d412, d413);
	buf ( d437, d41);
	nor ( d438, d410, d429);
	xor ( d439, d421, d427);
	nor ( d440, d411, d425);
	or ( d441, d416, d421);
	xor ( d442, d413, d429);
	nor ( d443, d411, d423);
	buf ( d444, d130);
	or ( d445, d420, d426);
	buf ( d446, d257);
	nand ( d447, d417, d424);
	xor ( d448, d417, d421);
	and ( d449, d418, d424);
	buf ( d450, d125);
	xor ( d451, d414, d415);
	not ( d452, d165);
	and ( d453, d413, d414);
	nor ( d454, d432, d444);
	nor ( d455, d434, d438);
	buf ( d456, d89);
	and ( d457, d434, d449);
	xnor ( d458, d444, d449);
	buf ( d459, d45);
	or ( d460, d445, d448);
	buf ( d461, d245);
	xnor ( d462, d433, d448);
	not ( d463, d330);
	or ( d464, d433, d439);
	xor ( d465, d435, d440);
	not ( d466, d439);
	xor ( d467, d461);
	and ( d468, d456, d458);
	nor ( d469, d459, d465);
	and ( d470, d459, d463);
	buf ( d471, d217);
	nand ( d472, d462, d464);
	nor ( d473, d457, d461);
	buf ( d474, d409);
	nor ( d475, d456, d463);
	not ( d476, d403);
	xor ( d477, d464);
	xnor ( d478, d454, d462);
	and ( d479, d455, d462);
	nand ( d480, d462, d465);
	nand ( d481, d460, d464);
	or ( d482, d454, d461);
	and ( d483, d455, d456);
	and ( d484, d455);
	xnor ( d485, d455, d456);
	nand ( d486, d463, d464);
	nor ( d487, d456, d465);
	or ( d488, d457);
	xor ( d489, d461, d462);
	and ( d490, d460, d464);
	nor ( d491, d459, d460);
	buf ( d492, d210);
	nor ( d493, d454, d464);
	not ( d494, d132);
	xnor ( d495, d457);
	xnor ( d496, d454);
	buf ( d497, d231);
	xnor ( d498, d461, d462);
	buf ( d499, d393);
	xor ( d500, d459, d461);
	not ( d501, d76);
	xor ( d502, d454, d463);
	or ( d503, d455, d459);
	not ( d504, d24);
	nand ( d505, d461, d464);
	nor ( d506, d456, d458);
	and ( d507, d457, d462);
	nand ( d508, d455, d457);
	or ( d509, d455, d461);
	or ( d510, d454, d455);
	xnor ( d511, d457, d462);
	xor ( d512, d455, d463);
	nand ( d513, d454, d457);
	buf ( d514, d5);
	xnor ( d515, d471, d492);
	and ( d516, d494, d510);
	xor ( d517, d474, d482);
	buf ( d518, d415);
	nand ( d519, d480, d489);
	and ( d520, d473, d485);
	or ( d521, d483, d503);
	nand ( d522, d471, d495);
	and ( d523, d477, d491);
	xnor ( d524, d482, d507);
	nand ( d525, d497, d508);
	xor ( d526, d471, d507);
	and ( d527, d471, d497);
	xor ( d528, d510, d511);
	not ( d529, d391);
	or ( d530, d481, d499);
	nand ( d531, d475, d476);
	xor ( d532, d466, d494);
	xnor ( d533, d472, d479);
	nor ( d534, d478, d483);
	nor ( d535, d466, d470);
	nand ( d536, d479, d496);
	xor ( d537, d487, d500);
	and ( d538, d467, d513);
	buf ( d539, d467);
	buf ( d540, d301);
	and ( d541, d466, d480);
	or ( d542, d471, d485);
	or ( d543, d478, d490);
	nand ( d544, d485, d505);
	or ( d545, d469, d504);
	or ( d546, d482, d488);
	xnor ( d547, d492, d500);
	buf ( d548, d484);
	or ( d549, d475, d494);
	not ( d550, d62);
	buf ( d551, d344);
	or ( d552, d489, d506);
	not ( d553, d459);
	nor ( d554, d471, d486);
	nand ( d555, d477, d499);
	nor ( d556, d468, d492);
	and ( d557, d472, d510);
	nor ( d558, d477, d481);
	nor ( d559, d471, d487);
	nand ( d560, d548, d559);
	nand ( d561, d556);
	not ( d562, d382);
	xnor ( d563, d546);
	nor ( d564, d533, d547);
	and ( d565, d522, d523);
	buf ( d566, d557);
	not ( d567, d11);
	not ( d568, d336);
	nand ( d569, d525, d528);
	or ( d570, d518, d538);
	nand ( d571, d521, d552);
	xnor ( d572, d542, d547);
	and ( d573, d520, d555);
	xnor ( d574, d569, d571);
	or ( d575, d565, d566);
	xnor ( d576, d561, d568);
	not ( d577, d437);
	or ( d578, d566);
	nand ( d579, d560, d570);
	xor ( d580, d576, d577);
	nand ( d581, d574);
	xor ( d582, d578, d579);
	xor ( d583, d577, d579);
	and ( d584, d575, d579);
	or ( d585, d577, d579);
	and ( d586, d576, d577);
	or ( d587, d575, d577);
	nand ( d588, d576, d577);
	buf ( d589, d252);
	buf ( d590, d401);
	xor ( d591, d575, d577);
	nor ( d592, d577, d578);
	not ( d593, d333);
	nor ( d594, d574, d575);
	nor ( d595, d577);
	nand ( d596, d575, d577);
	buf ( d597, d95);
	buf ( d598, d385);
	nand ( d599, d578, d579);
	not ( d600, d448);
	buf ( d601, d189);
	buf ( d602, d573);
	and ( d603, d587, d601);
	not ( d604, d226);
	buf ( d605, d330);
	nand ( d606, d583, d587);
	and ( d607, d585, d600);
	xor ( d608, d587, d592);
	or ( d609, d582, d602);
	xnor ( d610, d581);
	nor ( d611, d599, d601);
	xnor ( d612, d581, d590);
	or ( d613, d598, d602);
	buf ( d614, d542);
	or ( d615, d584, d601);
	xnor ( d616, d588, d600);
	not ( d617, d53);
	or ( d618, d591, d599);
	xnor ( d619, d589, d595);
	buf ( d620, d536);
	or ( d621, d590);
	and ( d622, d590, d602);
	buf ( d623, d357);
	not ( d624, d545);
	xnor ( d625, d590, d598);
	xnor ( d626, d587, d600);
	xnor ( d627, d582, d597);
	nand ( d628, d583, d593);
	nand ( d629, d582, d589);
	xor ( d630, d595, d598);
	or ( d631, d593, d597);
	xnor ( d632, d594, d602);
	buf ( d633, d60);
	nand ( d634, d591, d593);
	buf ( d635, d318);
	and ( d636, d581, d582);
	and ( d637, d582, d593);
	or ( d638, d594, d595);
	nand ( d639, d592, d595);
	xor ( d640, d580, d581);
	xnor ( d641, d586, d599);
	or ( d642, d597, d600);
	nor ( d643, d588, d589);
	nand ( d644, d586, d600);
	or ( d645, d585, d595);
	nor ( d646, d590);
	xnor ( d647, d591, d600);
	not ( d648, d35);
	xor ( d649, d608, d615);
	xnor ( d650, d625, d634);
	nand ( d651, d616, d630);
	xor ( d652, d609, d631);
	buf ( d653, d105);
	or ( d654, d605, d628);
	nand ( d655, d632, d636);
	and ( d656, d606, d614);
	buf ( d657, d203);
	or ( d658, d605, d626);
	or ( d659, d620, d646);
	and ( d660, d620, d632);
	and ( d661, d623, d624);
	xnor ( d662, d620, d642);
	nand ( d663, d638, d645);
	xor ( d664, d616, d631);
	buf ( d665, d516);
	nand ( d666, d624, d646);
	nand ( d667, d613, d642);
	or ( d668, d613, d619);
	not ( d669, d230);
	xnor ( d670, d611, d614);
	nand ( d671, d625, d630);
	nand ( d672, d621, d626);
	xor ( d673, d661, d664);
	nor ( d674, d648, d656);
	buf ( d675, d454);
	or ( d676, d655, d663);
	not ( d677, d369);
	xor ( d678, d650, d653);
	nand ( d679, d662, d670);
	or ( d680, d660, d670);
	nand ( d681, d648, d662);
	nor ( d682, d654, d671);
	buf ( d683, d55);
	nor ( d684, d658, d661);
	nor ( d685, d656, d666);
	or ( d686, d649, d658);
	and ( d687, d651, d656);
	nand ( d688, d650, d664);
	nand ( d689, d654, d666);
	xnor ( d690, d652, d655);
	nor ( d691, d658, d666);
	nor ( d692, d665, d668);
	xor ( d693, d650, d666);
	xnor ( d694, d660, d667);
	nor ( d695, d657, d662);
	or ( d696, d649, d650);
	and ( d697, d649, d662);
	xnor ( d698, d648, d661);
	xnor ( d699, d648, d670);
	xor ( d700, d661, d663);
	buf ( d701, d411);
	xnor ( d702, d661, d672);
	and ( d703, d662, d669);
	and ( d704, d662, d671);
	buf ( d705, d8);
	or ( d706, d665, d667);
	nor ( d707, d655, d670);
	xnor ( d708, d667, d672);
	nand ( d709, d661);
	and ( d710, d654, d657);
	not ( d711, d571);
	nand ( d712, d654, d666);
	nor ( d713, d665, d672);
	nand ( d714, d678, d689);
	nor ( d715, d674, d678);
	nand ( d716, d706, d708);
	nand ( d717, d680, d692);
	nand ( d718, d689, d693);
	nand ( d719, d700, d712);
	xor ( d720, d694, d698);
	nor ( d721, d681, d710);
	buf ( d722, d712);
	not ( d723, d171);
	nand ( d724, d680, d693);
	nor ( d725, d679, d686);
	nand ( d726, d689, d699);
	and ( d727, d675, d689);
	nand ( d728, d692, d694);
	not ( d729, d190);
	or ( d730, d694, d695);
	not ( d731, d205);
	buf ( d732, d541);
	nor ( d733, d674, d690);
	xor ( d734, d689);
	xnor ( d735, d702, d706);
	nor ( d736, d683, d685);
	xor ( d737, d681, d709);
	buf ( d738, d90);
	or ( d739, d691, d692);
	or ( d740, d692, d702);
	xnor ( d741, d688, d706);
	or ( d742, d702, d713);
	not ( d743, d700);
	nand ( d744, d673, d681);
	xnor ( d745, d686, d688);
	or ( d746, d683, d688);
	and ( d747, d677, d680);
	xnor ( d748, d687, d700);
	xnor ( d749, d694, d706);
	buf ( d750, d87);
	nor ( d751, d685, d690);
	not ( d752, d39);
	and ( d753, d698, d699);
	or ( d754, d674, d681);
	buf ( d755, d418);
	buf ( d756, d529);
	or ( d757, d724, d736);
	xnor ( d758, d729, d732);
	buf ( d759, d137);
	nand ( d760, d723, d736);
	xor ( d761, d715, d749);
	or ( d762, d729, d746);
	xnor ( d763, d733, d756);
	nor ( d764, d723, d749);
	xor ( d765, d732, d747);
	xnor ( d766, d730, d743);
	nand ( d767, d735, d752);
	xor ( d768, d737, d754);
	not ( d769, d564);
	buf ( d770, d632);
	xor ( d771, d720, d731);
	buf ( d772, d221);
	not ( d773, d449);
	not ( d774, d258);
	buf ( d775, d489);
	and ( d776, d714, d716);
	not ( d777, d678);
	nor ( d778, d717, d733);
	and ( d779, d716, d737);
	buf ( d780, d569);
	or ( d781, d725, d742);
	xnor ( d782, d728, d740);
	or ( d783, d735, d736);
	nor ( d784, d718, d732);
	nand ( d785, d725, d742);
	and ( d786, d714, d731);
	and ( d787, d770, d773);
	not ( d788, d358);
	not ( d789, d309);
	xor ( d790, d771, d786);
	nor ( d791, d763, d783);
	and ( d792, d760, d776);
	buf ( d793, d54);
	not ( d794, d51);
	not ( d795, d79);
	not ( d796, d48);
	nand ( d797, d772, d781);
	xnor ( d798, d774, d783);
	nand ( d799, d773, d774);
	xnor ( d800, d790, d794);
	nand ( d801, d789, d794);
	and ( d802, d789, d792);
	xnor ( d803, d797);
	xor ( d804, d798);
	or ( d805, d787, d793);
	xor ( d806, d789, d798);
	xnor ( d807, d793, d797);
	nand ( d808, d790);
	and ( d809, d798, d799);
	or ( d810, d791);
	and ( d811, d792, d797);
	nor ( d812, d792, d793);
	nor ( d813, d795, d797);
	buf ( d814, d229);
	xor ( d815, d792, d796);
	xnor ( d816, d790, d792);
	nand ( d817, d793, d799);
	or ( d818, d791, d799);
	or ( d819, d793, d799);
	buf ( d820, d795);
	xnor ( d821, d797, d798);
	not ( d822, d387);
	or ( d823, d794, d799);
	and ( d824, d795, d799);
	or ( d825, d789, d793);
	or ( d826, d789, d799);
	nor ( d827, d789, d792);
	nand ( d828, d788, d794);
	buf ( d829, d438);
	or ( d830, d794, d795);
	or ( d831, d791, d796);
	or ( d832, d789, d793);
	buf ( d833, d312);
	xnor ( d834, d791, d794);
	xor ( d835, d788, d789);
	assign f1 = d822;
	assign f2 = d825;
	assign f3 = d819;
	assign f4 = d820;
	assign f5 = d834;
	assign f6 = d818;
	assign f7 = d835;
	assign f8 = d810;
	assign f9 = d829;
	assign f10 = d813;
	assign f11 = d804;
	assign f12 = d823;
endmodule
