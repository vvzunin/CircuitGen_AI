module CCGRCG110( x0, x1, x2, x3, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17, f18, f19 );

	input x0, x1, x2, x3;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17, f18, f19;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314, d315, d316, d317, d318, d319, d320, d321, d322, d323, d324, d325, d326, d327, d328, d329, d330, d331, d332, d333, d334, d335, d336, d337, d338, d339, d340, d341, d342, d343, d344, d345, d346, d347, d348, d349, d350, d351, d352, d353, d354, d355, d356, d357, d358, d359, d360, d361, d362, d363, d364, d365, d366, d367, d368, d369, d370, d371, d372, d373, d374, d375, d376, d377, d378, d379, d380, d381, d382, d383, d384, d385, d386, d387, d388, d389, d390, d391, d392, d393, d394, d395, d396, d397, d398, d399, d400, d401, d402, d403, d404, d405, d406, d407, d408, d409, d410, d411, d412, d413, d414, d415, d416, d417, d418, d419, d420, d421, d422, d423, d424, d425, d426, d427, d428, d429, d430, d431, d432, d433, d434, d435, d436, d437, d438, d439, d440, d441, d442, d443, d444, d445, d446, d447, d448, d449, d450, d451;

	xor (d1, x0, x3);
	nor (d2, x0, x1);
	nand (d3, x0, x1);
	buf (d4, x3);
	nand (d5, x2, x3);
	xor (d6, x0);
	not (d7, x2);
	or (d8, x0, x3);
	or (d9, x0, x3);
	xor (d10, x1, x3);
	nor (d11, x3);
	nor (d12, x2, x3);
	or (d13, x1, x3);
	nand (d14, x1);
	and (d15, x1, x3);
	buf (d16, x1);
	and (d17, x1, x3);
	xnor (d18, x1);
	xnor (d19, x1, x3);
	xnor (d20, x2);
	not (d21, x1);
	xor (d22, x0, x2);
	xor (d23, x2);
	xor (d24, x0, x3);
	or (d25, x0, x2);
	nand (d26, x1, x3);
	not (d27, x3);
	xor (d28, d14, d26);
	buf (d29, d18);
	or (d30, d7, d25);
	or (d31, d16);
	xor (d32, d11, d20);
	not (d33, d4);
	buf (d34, d19);
	not (d35, d8);
	xor (d36, d4, d26);
	not (d37, d15);
	nand (d38, d5, d18);
	xnor (d39, d3, d18);
	or (d40, d6, d26);
	xnor (d41, d13, d17);
	nand (d42, d1, d3);
	nand (d43, d2, d5);
	nand (d44, d6, d27);
	xor (d45, d7, d13);
	or (d46, d7, d16);
	or (d47, d2, d6);
	not (d48, d19);
	nor (d49, d13, d19);
	or (d50, d6, d27);
	not (d51, d24);
	nand (d52, d1, d7);
	buf (d53, d9);
	xnor (d54, d3, d7);
	xor (d55, d3, d5);
	and (d56, d15, d20);
	nor (d57, d12, d25);
	buf (d58, d6);
	or (d59, d23);
	not (d60, d3);
	xor (d61, d4, d23);
	nor (d62, d9, d16);
	xnor (d63, d3, d13);
	and (d64, d17, d22);
	and (d65, d14, d17);
	nor (d66, d19, d22);
	buf (d67, d24);
	xnor (d68, d3, d8);
	nor (d69, d8, d10);
	or (d70, d1, d26);
	nor (d71, d9, d18);
	xnor (d72, d19, d20);
	nor (d73, d3, d20);
	xnor (d74, d6, d18);
	nand (d75, d7, d23);
	and (d76, d4, d17);
	and (d77, d1, d17);
	xor (d78, d12, d18);
	or (d79, d1, d12);
	buf (d80, d16);
	or (d81, d7, d12);
	and (d82, d14, d23);
	xor (d83, d3, d27);
	or (d84, d20, d22);
	nor (d85, d3, d16);
	buf (d86, d15);
	not (d87, d48);
	and (d88, d48, d78);
	not (d89, d85);
	xor (d90, d61, d70);
	nand (d91, d33, d83);
	nand (d92, d37, d69);
	nand (d93, d53, d80);
	nand (d94, d64, d81);
	not (d95, d14);
	xor (d96, d80);
	xor (d97, d62, d79);
	xor (d98, d34, d52);
	xor (d99, d43, d68);
	nor (d100, d32, d57);
	not (d101, d57);
	xnor (d102, d46, d73);
	xnor (d103, d50, d65);
	not (d104, d9);
	nand (d105, d30, d33);
	and (d106, d46, d64);
	and (d107, d51, d71);
	and (d108, d58, d64);
	buf (d109, d29);
	xor (d110, d63, d80);
	xor (d111, d57, d85);
	buf (d112, d14);
	xnor (d113, d59, d79);
	nor (d114, d30, d59);
	xor (d115, d37, d72);
	xor (d116, d46, d49);
	nand (d117, d34, d74);
	xor (d118, d61, d76);
	not (d119, d33);
	nor (d120, d34, d60);
	nand (d121, d61, d86);
	or (d122, d58, d64);
	not (d123, d36);
	or (d124, d52, d60);
	and (d125, d35, d51);
	or (d126, d69, d75);
	and (d127, d47, d65);
	nand (d128, d43, d84);
	not (d129, d39);
	xor (d130, d41, d63);
	and (d131, d80, d85);
	buf (d132, d43);
	or (d133, d39, d71);
	not (d134, d50);
	xor (d135, d39, d75);
	buf (d136, d85);
	buf (d137, d50);
	and (d138, d38, d74);
	xor (d139, d67, d86);
	xnor (d140, d33, d76);
	xor (d141, d73, d76);
	buf (d142, d35);
	nor (d143, d40, d53);
	not (d144, d16);
	buf (d145, d60);
	buf (d146, d86);
	xnor (d147, d49, d53);
	nand (d148, d46, d66);
	buf (d149, d41);
	nand (d150, d76, d85);
	not (d151, d86);
	not (d152, d72);
	nand (d153, d32, d58);
	xnor (d154, d45, d51);
	nand (d155, d41, d75);
	nand (d156, d37, d45);
	or (d157, d29, d48);
	xor (d158, d51, d57);
	or (d159, d51, d76);
	not (d160, d26);
	nand (d161, d149, d152);
	nand (d162, d121, d141);
	not (d163, d102);
	nand (d164, d97, d159);
	or (d165, d102, d128);
	or (d166, d92, d114);
	nor (d167, d99, d144);
	xor (d168, d122, d139);
	nand (d169, d92, d130);
	buf (d170, d67);
	nand (d171, d99, d104);
	or (d172, d121, d155);
	xnor (d173, d104, d144);
	nand (d174, d88, d104);
	not (d175, d154);
	not (d176, d42);
	or (d177, d138, d142);
	xor (d178, d100, d139);
	and (d179, d110, d136);
	not (d180, d160);
	not (d181, d145);
	not (d182, d28);
	not (d183, d56);
	and (d184, d91, d108);
	or (d185, d99, d141);
	xor (d186, d138, d140);
	xor (d187, d124, d131);
	nand (d188, d145, d159);
	buf (d189, d53);
	buf (d190, d146);
	nor (d191, d97, d134);
	buf (d192, d154);
	or (d193, d110, d143);
	or (d194, d110, d136);
	and (d195, d112, d117);
	xnor (d196, d149, d158);
	nor (d197, d94, d117);
	not (d198, d75);
	or (d199, d137, d148);
	buf (d200, d96);
	and (d201, d105, d143);
	nor (d202, d108, d129);
	nor (d203, d104, d153);
	or (d204, d107, d148);
	and (d205, d122, d135);
	xor (d206, d129, d151);
	nor (d207, d104, d128);
	xnor (d208, d97, d142);
	buf (d209, d160);
	xor (d210, d101, d121);
	xnor (d211, d92, d141);
	xnor (d212, d125, d157);
	not (d213, d112);
	not (d214, d11);
	xnor (d215, d110, d154);
	xnor (d216, d162, d174);
	nand (d217, d168, d202);
	xnor (d218, d179, d186);
	buf (d219, d202);
	not (d220, d129);
	buf (d221, d139);
	buf (d222, d77);
	xnor (d223, d164, d168);
	nor (d224, d179, d203);
	or (d225, d183, d207);
	nand (d226, d171, d214);
	not (d227, d139);
	or (d228, d163, d190);
	nand (d229, d195, d214);
	xnor (d230, d161, d172);
	buf (d231, d125);
	xnor (d232, d168, d206);
	nand (d233, d179, d187);
	xor (d234, d181, d194);
	nor (d235, d186, d200);
	xnor (d236, d178, d211);
	xor (d237, d176, d189);
	xor (d238, d179);
	and (d239, d201, d208);
	nor (d240, d181, d211);
	not (d241, d95);
	buf (d242, d57);
	nand (d243, d168, d183);
	xnor (d244, d198);
	buf (d245, d192);
	and (d246, d179, d202);
	nand (d247, d178, d213);
	xor (d248, d219, d220);
	and (d249, d218, d247);
	and (d250, d222, d233);
	xor (d251, d220, d226);
	nor (d252, d225, d229);
	xor (d253, d229, d232);
	buf (d254, d230);
	nor (d255, d225, d234);
	buf (d256, d194);
	nor (d257, d233, d240);
	xnor (d258, d227, d238);
	not (d259, d247);
	xnor (d260, d236, d242);
	buf (d261, d7);
	nor (d262, d225, d238);
	nor (d263, d234, d235);
	nand (d264, d216, d231);
	xor (d265, d224, d242);
	nand (d266, d221, d245);
	not (d267, d108);
	nor (d268, d230, d246);
	xor (d269, d217, d236);
	buf (d270, d195);
	nor (d271, d241, d244);
	nor (d272, d224, d226);
	buf (d273, d100);
	not (d274, d203);
	and (d275, d232, d238);
	xor (d276, d217, d221);
	xor (d277, d219, d237);
	nor (d278, d220, d245);
	nor (d279, d218, d232);
	and (d280, d227, d237);
	not (d281, d201);
	xnor (d282, d221, d224);
	nor (d283, d224, d247);
	nand (d284, d219, d224);
	or (d285, d220, d229);
	nor (d286, d224, d232);
	buf (d287, d144);
	not (d288, d103);
	nand (d289, d222, d245);
	xor (d290, d219, d239);
	nor (d291, d242, d247);
	xnor (d292, d225, d246);
	nand (d293, d243, d246);
	and (d294, d220, d246);
	xnor (d295, d218, d240);
	or (d296, d219, d225);
	nand (d297, d226, d244);
	not (d298, d148);
	buf (d299, d113);
	nor (d300, d217, d244);
	nor (d301, d220, d225);
	not (d302, d99);
	nand (d303, d241, d243);
	xnor (d304, d223, d233);
	or (d305, d222, d223);
	xnor (d306, d241, d246);
	not (d307, d230);
	nor (d308, d230, d240);
	xor (d309, d241, d245);
	or (d310, d227, d233);
	buf (d311, d111);
	nand (d312, d216, d237);
	nand (d313, d226, d232);
	or (d314, d216, d244);
	or (d315, d226, d246);
	nor (d316, d232, d238);
	or (d317, d227, d234);
	nand (d318, d220, d226);
	nand (d319, d220, d234);
	or (d320, d231, d242);
	buf (d321, d157);
	buf (d322, d215);
	or (d323, d217, d244);
	not (d324, d207);
	nor (d325, d216, d246);
	nand (d326, d221, d224);
	not (d327, d43);
	xor (d328, d236, d243);
	nand (d329, d217, d246);
	buf (d330, d203);
	and (d331, d217, d240);
	nor (d332, d270, d304);
	nand (d333, d250, d322);
	and (d334, d308, d324);
	nor (d335, d274, d312);
	xnor (d336, d305, d323);
	xor (d337, d264, d323);
	nor (d338, d255, d328);
	nor (d339, d264, d291);
	and (d340, d261, d280);
	nand (d341, d283, d316);
	or (d342, d299, d319);
	nor (d343, d308, d319);
	not (d344, d93);
	nand (d345, d313);
	not (d346, d240);
	xnor (d347, d268, d282);
	and (d348, d251, d320);
	xnor (d349, d269, d292);
	nor (d350, d292, d331);
	or (d351, d303, d320);
	or (d352, d280, d284);
	xor (d353, d300, d318);
	or (d354, d273, d290);
	xnor (d355, d253, d316);
	nand (d356, d261, d279);
	and (d357, d280, d307);
	buf (d358, d132);
	xnor (d359, d344, d349);
	and (d360, d347, d348);
	or (d361, d347, d352);
	xnor (d362, d334, d335);
	xnor (d363, d347, d349);
	or (d364, d333, d347);
	and (d365, d344, d349);
	nor (d366, d345, d350);
	not (d367, d146);
	or (d368, d337, d349);
	buf (d369, d265);
	nand (d370, d342, d351);
	and (d371, d339, d348);
	not (d372, d325);
	or (d373, d333, d343);
	nor (d374, d350, d357);
	nor (d375, d333, d341);
	nand (d376, d337, d354);
	xnor (d377, d340, d355);
	not (d378, d209);
	buf (d379, d78);
	buf (d380, d131);
	and (d381, d337, d351);
	or (d382, d333, d349);
	buf (d383, d180);
	and (d384, d338, d342);
	nand (d385, d333, d346);
	or (d386, d336, d349);
	buf (d387, d232);
	or (d388, d346, d351);
	buf (d389, d115);
	xnor (d390, d343, d345);
	nor (d391, d345, d346);
	or (d392, d341, d350);
	xor (d393, d346, d351);
	buf (d394, d22);
	xnor (d395, d348);
	nor (d396, d342, d350);
	xnor (d397, d352, d356);
	xnor (d398, d338, d340);
	or (d399, d344, d352);
	nand (d400, d334, d351);
	xor (d401, d333, d345);
	nor (d402, d345, d347);
	nand (d403, d353, d354);
	and (d404, d355, d356);
	buf (d405, d267);
	buf (d406, d109);
	nand (d407, d340, d347);
	xor (d408, d347, d352);
	and (d409, d351, d356);
	and (d410, d337, d357);
	and (d411, d357);
	xor (d412, d336, d357);
	nor (d413, d349, d356);
	nor (d414, d332, d337);
	nor (d415, d355, d356);
	xnor (d416, d340, d351);
	nand (d417, d336, d339);
	and (d418, d341, d346);
	nand (d419, d336, d346);
	not (d420, d327);
	buf (d421, d142);
	xnor (d422, d343, d353);
	xnor (d423, d335, d342);
	and (d424, d333, d339);
	xor (d425, d352, d356);
	nand (d426, d340, d355);
	or (d427, d334, d335);
	xnor (d428, d333, d344);
	and (d429, d349, d354);
	xnor (d430, d333, d355);
	not (d431, d274);
	xnor (d432, d339, d352);
	xor (d433, d342, d355);
	buf (d434, d20);
	nand (d435, d337, d356);
	buf (d436, d283);
	and (d437, d344, d354);
	xor (d438, d334, d350);
	and (d439, d340, d351);
	xor (d440, d337, d357);
	xor (d441, d343, d352);
	or (d442, d336, d356);
	or (d443, d336, d339);
	xnor (d444, d337, d345);
	xor (d445, d343, d347);
	and (d446, d333, d346);
	not (d447, d295);
	xnor (d448, d333, d354);
	xor (d449, d338, d357);
	nor (d450, d337, d347);
	nor (d451, d341, d350);
	assign f1 = d448;
	assign f2 = d413;
	assign f3 = d381;
	assign f4 = d373;
	assign f5 = d435;
	assign f6 = d440;
	assign f7 = d430;
	assign f8 = d393;
	assign f9 = d417;
	assign f10 = d373;
	assign f11 = d374;
	assign f12 = d404;
	assign f13 = d434;
	assign f14 = d392;
	assign f15 = d384;
	assign f16 = d363;
	assign f17 = d390;
	assign f18 = d416;
	assign f19 = d432;
endmodule
