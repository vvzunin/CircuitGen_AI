module CCGRCG95( x0, x1, x2, x3, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11 );

	input x0, x1, x2, x3;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314, d315, d316, d317, d318, d319, d320, d321, d322, d323, d324, d325, d326, d327, d328, d329, d330, d331, d332, d333, d334, d335, d336, d337, d338, d339, d340, d341, d342, d343, d344, d345, d346, d347, d348, d349, d350, d351, d352, d353, d354, d355, d356, d357, d358, d359, d360, d361, d362, d363, d364, d365, d366, d367, d368, d369, d370, d371, d372, d373, d374, d375, d376, d377, d378, d379, d380, d381, d382, d383, d384, d385, d386, d387, d388, d389, d390, d391, d392, d393, d394, d395, d396, d397, d398, d399, d400, d401, d402, d403, d404, d405, d406, d407, d408, d409, d410, d411, d412, d413, d414, d415, d416, d417, d418, d419, d420, d421, d422, d423, d424, d425, d426, d427, d428, d429, d430, d431, d432, d433, d434, d435, d436, d437, d438, d439, d440, d441, d442, d443, d444, d445, d446, d447, d448, d449, d450, d451, d452, d453, d454, d455, d456, d457, d458, d459, d460, d461, d462, d463, d464, d465, d466, d467, d468, d469, d470, d471, d472, d473, d474, d475, d476, d477, d478, d479, d480, d481, d482, d483, d484, d485, d486, d487, d488, d489, d490, d491, d492, d493, d494, d495, d496, d497, d498, d499, d500, d501, d502, d503, d504;

	or (d1, x0, x3);
	not (d2, x3);
	buf (d3, x3);
	or (d4, x1);
	or (d5, x1, x3);
	xor (d6, x1, x3);
	nor (d7, x1, x2);
	not (d8, x0);
	nand (d9, x1);
	nor (d10, x0, x2);
	and (d11, x0, x3);
	or (d12, x2);
	xnor (d13, x0, x2);
	nor (d14, x2, x3);
	nand (d15, x1, x3);
	nand (d16, x0, x1);
	xnor (d17, x1);
	xnor (d18, x0);
	nand (d19, x2, x3);
	nand (d20, x3);
	or (d21, x0, x1);
	nand (d22, d1);
	not (d23, d19);
	xor (d24, d8, d13);
	nor (d25, d8, d21);
	xnor (d26, d6, d12);
	xnor (d27, d8, d19);
	not (d28, d9);
	nand (d29, d19, d20);
	nor (d30, d5, d11);
	buf (d31, x0);
	and (d32, d11, d19);
	xor (d33, d4, d16);
	nand (d34, d14, d18);
	not (d35, d8);
	xnor (d36, d1, d3);
	nor (d37, d1, d19);
	and (d38, d9, d14);
	buf (d39, d2);
	nand (d40, d7, d11);
	or (d41, d25, d40);
	xnor (d42, d34, d38);
	or (d43, d24, d27);
	nor (d44, d24, d39);
	nand (d45, d24, d36);
	xnor (d46, d24, d30);
	xor (d47, d26, d27);
	xor (d48, d31, d35);
	nand (d49, d27, d31);
	and (d50, d22, d35);
	xnor (d51, d35, d38);
	not (d52, d39);
	xnor (d53, d23, d36);
	buf (d54, d32);
	xnor (d55, d34, d37);
	nor (d56, d22, d35);
	xnor (d57, d22, d38);
	nor (d58, d29, d40);
	xor (d59, d31, d33);
	or (d60, d33, d39);
	nand (d61, d36, d39);
	or (d62, d24, d38);
	nor (d63, d26, d39);
	nand (d64, d31, d32);
	nor (d65, d32, d38);
	nand (d66, d32, d35);
	nand (d67, d23, d30);
	buf (d68, d38);
	buf (d69, d29);
	nor (d70, d26, d27);
	nor (d71, d25, d29);
	xor (d72, d25, d28);
	xor (d73, d28, d32);
	and (d74, d23, d36);
	buf (d75, d6);
	buf (d76, d37);
	and (d77, d27, d30);
	nor (d78, d31, d35);
	buf (d79, d18);
	xor (d80, d22);
	and (d81, d26, d38);
	xnor (d82, d22, d38);
	buf (d83, d23);
	nand (d84, d33, d39);
	xor (d85, d25, d39);
	or (d86, d30, d40);
	not (d87, d36);
	xor (d88, d47, d84);
	or (d89, d51, d71);
	buf (d90, d25);
	xor (d91, d62, d65);
	or (d92, d53, d83);
	nand (d93, d41, d44);
	xnor (d94, d61, d66);
	or (d95, d67, d83);
	xor (d96, d69, d74);
	nand (d97, d61, d62);
	xnor (d98, d47, d73);
	nand (d99, d72, d77);
	buf (d100, d28);
	and (d101, d63, d73);
	xor (d102, d41, d45);
	nor (d103, d46, d66);
	nor (d104, d64, d85);
	nand (d105, d53, d80);
	nor (d106, d63, d73);
	or (d107, d49, d66);
	and (d108, d53, d77);
	nand (d109, d46, d71);
	or (d110, d77, d84);
	not (d111, d82);
	not (d112, d55);
	nor (d113, d58, d70);
	or (d114, d59);
	nand (d115, d43, d49);
	nand (d116, d69, d76);
	nand (d117, d50, d68);
	xor (d118, d70, d75);
	nand (d119, d57, d81);
	xor (d120, d75, d83);
	not (d121, d35);
	xnor (d122, d53, d86);
	xnor (d123, d62, d68);
	nand (d124, d44, d46);
	nand (d125, d67, d86);
	nor (d126, d60, d85);
	or (d127, d58, d70);
	or (d128, d71, d78);
	buf (d129, d19);
	nand (d130, d52, d65);
	and (d131, d47, d63);
	nand (d132, d49, d81);
	xor (d133, d47, d57);
	and (d134, d60, d81);
	and (d135, d102, d115);
	nor (d136, d118, d130);
	and (d137, d113, d120);
	nand (d138, d103, d109);
	and (d139, d87, d133);
	buf (d140, d132);
	not (d141, d117);
	or (d142, d105, d114);
	and (d143, d93, d114);
	or (d144, d97, d123);
	xnor (d145, d107, d121);
	buf (d146, d10);
	and (d147, d113, d118);
	xor (d148, d87, d99);
	xnor (d149, d112, d129);
	xor (d150, d88, d113);
	or (d151, d112, d123);
	not (d152, d45);
	nand (d153, d102, d109);
	xor (d154, d122, d129);
	not (d155, d25);
	xor (d156, d94, d128);
	nand (d157, d98, d107);
	nor (d158, d98, d101);
	nor (d159, d120, d121);
	xnor (d160, d88, d133);
	nor (d161, d93, d112);
	xor (d162, d125, d127);
	buf (d163, d95);
	buf (d164, d12);
	and (d165, d121, d125);
	nor (d166, d93, d132);
	and (d167, d91, d124);
	and (d168, d124, d125);
	or (d169, d99, d126);
	xor (d170, d92, d101);
	not (d171, d64);
	nand (d172, d100, d109);
	nand (d173, d89, d103);
	xnor (d174, d108, d124);
	nor (d175, d102, d112);
	not (d176, d11);
	or (d177, d99, d103);
	nand (d178, d88, d93);
	and (d179, d101, d126);
	nand (d180, d137, d164);
	or (d181, d161, d173);
	xnor (d182, d161, d175);
	nand (d183, d141, d163);
	xnor (d184, d139, d159);
	nand (d185, d150, d163);
	buf (d186, d53);
	or (d187, d165, d172);
	and (d188, d150, d167);
	and (d189, d162, d176);
	not (d190, d50);
	nor (d191, d139, d146);
	nor (d192, d138, d154);
	buf (d193, d86);
	nor (d194, d137, d146);
	xor (d195, d149, d162);
	not (d196, d134);
	xnor (d197, d154, d165);
	buf (d198, d116);
	xor (d199, d137, d177);
	and (d200, d141, d161);
	buf (d201, d114);
	not (d202, d118);
	nand (d203, d157, d166);
	or (d204, d168, d170);
	and (d205, d141, d157);
	xor (d206, d142, d172);
	nand (d207, d157, d167);
	nand (d208, d136, d137);
	and (d209, d153, d167);
	and (d210, d151, d162);
	nand (d211, d139, d147);
	and (d212, d160, d179);
	nor (d213, d165, d176);
	xnor (d214, d151, d176);
	nor (d215, d143, d169);
	or (d216, d144, d155);
	xnor (d217, d140, d159);
	nor (d218, d135, d163);
	nor (d219, d191, d213);
	nand (d220, d216, d217);
	or (d221, d215, d218);
	xor (d222, d188, d217);
	xnor (d223, d196, d207);
	or (d224, d185, d205);
	xor (d225, d190, d213);
	xor (d226, d187, d215);
	nand (d227, d186, d207);
	buf (d228, d212);
	nand (d229, d208, d218);
	and (d230, d212);
	and (d231, d194);
	buf (d232, d101);
	nor (d233, d186, d212);
	nand (d234, d180, d202);
	xnor (d235, d199, d202);
	xnor (d236, d182, d187);
	nor (d237, d187, d197);
	buf (d238, d166);
	nor (d239, d190, d203);
	not (d240, d3);
	nand (d241, d199, d218);
	nor (d242, d197, d201);
	and (d243, d183, d202);
	not (d244, d108);
	nand (d245, d197, d206);
	nand (d246, d181, d195);
	and (d247, d209);
	or (d248, d192, d216);
	buf (d249, d211);
	nand (d250, d193, d213);
	nor (d251, d193, d213);
	nand (d252, d191, d204);
	xor (d253, d202, d212);
	nand (d254, d191, d207);
	not (d255, d6);
	buf (d256, d205);
	buf (d257, d64);
	buf (d258, d87);
	not (d259, d119);
	nor (d260, d186, d199);
	xor (d261, d189, d209);
	xor (d262, d181, d202);
	and (d263, d188, d199);
	xnor (d264, d203, d208);
	xnor (d265, d182, d202);
	not (d266, d89);
	nor (d267, d180, d206);
	not (d268, d57);
	not (d269, d139);
	or (d270, d195, d198);
	xnor (d271, d190, d215);
	not (d272, d80);
	not (d273, d70);
	buf (d274, d103);
	xnor (d275, d198, d215);
	nand (d276, d206, d216);
	xnor (d277, d183, d194);
	or (d278, d204, d215);
	xor (d279, d185, d199);
	xnor (d280, d183, d200);
	nor (d281, d206, d218);
	or (d282, d213, d217);
	xor (d283, d189, d190);
	xnor (d284, d204, d207);
	xor (d285, d193, d201);
	nor (d286, d204, d205);
	buf (d287, d147);
	xor (d288, d191, d218);
	nor (d289, d208, d216);
	and (d290, d181, d213);
	nor (d291, d186, d187);
	and (d292, d199, d210);
	not (d293, d187);
	or (d294, d184, d187);
	nor (d295, d183, d211);
	xor (d296, d203, d218);
	nor (d297, d206, d211);
	buf (d298, d161);
	xor (d299, d203, d208);
	xnor (d300, d189, d198);
	not (d301, d40);
	or (d302, d185, d197);
	not (d303, d65);
	not (d304, d163);
	and (d305, d211, d213);
	nand (d306, d211, d216);
	nor (d307, d200, d214);
	nor (d308, d195, d196);
	nor (d309, d211, d218);
	or (d310, d206, d207);
	xnor (d311, d214, d216);
	buf (d312, d56);
	buf (d313, d15);
	and (d314, d181, d183);
	xnor (d315, d180, d214);
	xor (d316, d180, d209);
	nand (d317, d231, d253);
	xnor (d318, d233, d289);
	xor (d319, d287, d307);
	and (d320, d219, d281);
	nand (d321, d238, d272);
	buf (d322, d62);
	and (d323, d251, d272);
	buf (d324, d168);
	nor (d325, d265, d300);
	not (d326, d212);
	nor (d327, d284, d301);
	nand (d328, d226, d283);
	or (d329, d221, d269);
	xnor (d330, d249, d254);
	xnor (d331, d241, d262);
	or (d332, d221, d285);
	or (d333, d289, d315);
	nand (d334, d219, d275);
	not (d335, d280);
	and (d336, d288, d308);
	not (d337, d170);
	xnor (d338, d286, d315);
	or (d339, d262, d299);
	not (d340, d254);
	nor (d341, d231, d281);
	nor (d342, d303, d316);
	buf (d343, d200);
	or (d344, d267, d268);
	or (d345, d219, d261);
	nand (d346, d242, d243);
	and (d347, d225, d272);
	xor (d348, d261, d298);
	xnor (d349, d292, d302);
	xor (d350, d238, d261);
	and (d351, d252, d274);
	buf (d352, d295);
	nor (d353, d277, d293);
	xor (d354, d301, d309);
	buf (d355, d100);
	or (d356, d226, d232);
	nor (d357, d245, d255);
	xor (d358, d281, d294);
	not (d359, d54);
	nand (d360, d260, d261);
	not (d361, d157);
	xor (d362, d258, d283);
	or (d363, d234, d246);
	not (d364, d111);
	and (d365, d274, d290);
	and (d366, d246, d277);
	nand (d367, d254, d299);
	nand (d368, d251, d311);
	xnor (d369, d222, d235);
	not (d370, d226);
	buf (d371, d140);
	or (d372, d247, d281);
	not (d373, d250);
	buf (d374, d156);
	not (d375, d110);
	or (d376, d261, d305);
	and (d377, d227, d232);
	nand (d378, d249, d259);
	xnor (d379, d238, d263);
	nand (d380, d245, d309);
	nand (d381, d286, d304);
	nor (d382, d351, d357);
	nor (d383, d357, d364);
	and (d384, d325);
	and (d385, d326, d357);
	and (d386, d320, d376);
	nor (d387, d333, d337);
	xnor (d388, d317, d346);
	or (d389, d322, d357);
	nand (d390, d336, d364);
	and (d391, d374, d376);
	not (d392, d217);
	buf (d393, d104);
	not (d394, d246);
	and (d395, d360, d375);
	xor (d396, d327, d360);
	not (d397, d281);
	xor (d398, d333, d380);
	xor (d399, d326, d350);
	or (d400, d334, d372);
	xnor (d401, d346, d369);
	not (d402, d84);
	not (d403, d41);
	xor (d404, d359, d380);
	nor (d405, d361, d363);
	nor (d406, d321, d368);
	nor (d407, d321, d356);
	and (d408, d351, d377);
	nand (d409, d323, d357);
	not (d410, d271);
	nand (d411, d328, d356);
	nor (d412, d319, d351);
	xor (d413, d368, d376);
	or (d414, d351, d355);
	nor (d415, d348, d366);
	nor (d416, d318, d379);
	and (d417, d339, d367);
	and (d418, d323, d335);
	nor (d419, d322, d351);
	nor (d420, d341, d346);
	nand (d421, d328, d347);
	xor (d422, d321, d345);
	or (d423, d360, d376);
	buf (d424, d24);
	xnor (d425, d341, d362);
	nand (d426, d347, d371);
	buf (d427, d194);
	nand (d428, d352, d371);
	nand (d429, d322, d341);
	xor (d430, d338, d378);
	nor (d431, d339, d364);
	nand (d432, d325, d356);
	not (d433, d161);
	buf (d434, d115);
	xnor (d435, d332, d333);
	or (d436, d335, d363);
	and (d437, d331, d345);
	nor (d438, d354, d377);
	nor (d439, d341, d359);
	not (d440, d366);
	xnor (d441, d333, d352);
	nor (d442, d351, d356);
	xnor (d443, d384, d441);
	and (d444, d425, d429);
	not (d445, x1);
	and (d446, d395, d414);
	and (d447, d417, d442);
	or (d448, d397, d430);
	nand (d449, d408, d435);
	not (d450, d93);
	xnor (d451, d395, d424);
	nor (d452, d408, d433);
	buf (d453, d403);
	or (d454, d401, d414);
	not (d455, d284);
	buf (d456, d294);
	nor (d457, d382, d442);
	not (d458, d356);
	buf (d459, d119);
	xnor (d460, d393, d426);
	nor (d461, d434, d438);
	xnor (d462, d383, d415);
	nand (d463, d401, d440);
	and (d464, d392, d395);
	xor (d465, d382, d389);
	nand (d466, d385, d405);
	not (d467, d426);
	not (d468, d240);
	and (d469, d390, d423);
	and (d470, d383, d387);
	and (d471, d403, d430);
	buf (d472, d371);
	not (d473, d438);
	buf (d474, d368);
	xor (d475, d384, d395);
	nor (d476, d394, d413);
	or (d477, d389, d438);
	and (d478, d412, d441);
	xnor (d479, d385, d402);
	xnor (d480, d398, d405);
	xnor (d481, d422);
	and (d482, d399, d428);
	not (d483, d154);
	or (d484, d392, d430);
	or (d485, d384, d430);
	or (d486, d384, d427);
	not (d487, d417);
	and (d488, d390, d431);
	and (d489, d384, d422);
	and (d490, d433, d437);
	xnor (d491, d405, d431);
	and (d492, d392, d425);
	not (d493, d346);
	xor (d494, d407, d416);
	and (d495, d434, d441);
	and (d496, d385, d416);
	nor (d497, d387, d395);
	xor (d498, d395, d410);
	xor (d499, d422, d423);
	nor (d500, d385, d427);
	not (d501, d435);
	nor (d502, d430, d435);
	xor (d503, d404, d436);
	and (d504, d423, d435);
	assign f1 = d486;
	assign f2 = d449;
	assign f3 = d490;
	assign f4 = d492;
	assign f5 = d469;
	assign f6 = d447;
	assign f7 = d473;
	assign f8 = d477;
	assign f9 = d443;
	assign f10 = d496;
	assign f11 = d461;
endmodule
