module CCGRCG97( x0, x1, x2, x3, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12 );

	input x0, x1, x2, x3;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157;

	buf (d1, x2);
	xnor (d2, x1, x3);
	and (d3, x0, x2);
	xor (d4, x1);
	nor (d5, x1, x2);
	xnor (d6, x2, x3);
	buf (d7, x0);
	nor (d8, x3);
	or (d9, x1, x3);
	not (d10, d9);
	nand (d11, d3);
	nor (d12, d4, d8);
	nor (d13, d2, d4);
	or (d14, d2, d4);
	nand (d15, d1, d2);
	nand (d16, d3, d7);
	xnor (d17, d2, d3);
	nand (d18, d12, d17);
	xnor (d19, d10, d12);
	or (d20, d11, d14);
	not (d21, d6);
	nand (d22, d15);
	buf (d23, d16);
	xnor (d24, d10, d11);
	or (d25, d12, d15);
	xor (d26, d11, d12);
	xnor (d27, d13, d16);
	xnor (d28, d15, d16);
	buf (d29, d13);
	xnor (d30, d13);
	nor (d31, d13, d17);
	xnor (d32, d13, d17);
	buf (d33, x1);
	xnor (d34, d15, d17);
	or (d35, d11, d13);
	not (d36, d5);
	and (d37, d15, d17);
	xor (d38, d11, d12);
	xor (d39, d15, d16);
	nand (d40, d13, d16);
	or (d41, d13, d14);
	and (d42, d13);
	nor (d43, d10, d14);
	not (d44, d1);
	not (d45, d3);
	nand (d46, d13, d15);
	buf (d47, d4);
	nand (d48, d11, d16);
	nand (d49, d13);
	and (d50, d10, d16);
	buf (d51, d1);
	and (d52, d14, d15);
	xor (d53, d10, d17);
	xor (d54, d12, d13);
	nand (d55, d10, d16);
	and (d56, d10);
	xnor (d57, d10);
	xnor (d58, d16, d17);
	nor (d59, d12, d17);
	xnor (d60, d15, d16);
	and (d61, d13, d17);
	nand (d62, d10, d16);
	xor (d63, d11, d17);
	or (d64, d10);
	xnor (d65, d11, d14);
	not (d66, x0);
	and (d67, d11, d14);
	or (d68, d15, d17);
	or (d69, d10, d11);
	nor (d70, d12);
	xor (d71, d13, d17);
	xnor (d72, d13, d14);
	buf (d73, d12);
	and (d74, d10, d11);
	xnor (d75, d16, d17);
	and (d76, d13, d15);
	xor (d77, d11, d15);
	or (d78, d15, d16);
	nand (d79, d12, d14);
	nand (d80, d10, d12);
	or (d81, d12, d14);
	buf (d82, d6);
	not (d83, d13);
	buf (d84, x3);
	not (d85, d12);
	xor (d86, d10, d16);
	nor (d87, d14, d16);
	not (d88, x3);
	or (d89, d12, d13);
	nor (d90, d10, d11);
	xnor (d91, d11, d16);
	nor (d92, d13);
	nor (d93, d11);
	buf (d94, d14);
	not (d95, x1);
	xnor (d96, d11, d17);
	nor (d97, d11, d15);
	not (d98, d2);
	nor (d99, d42, d52);
	and (d100, d64, d93);
	nand (d101, d43, d59);
	xor (d102, d32, d83);
	xor (d103, d57, d70);
	or (d104, d31, d85);
	and (d105, d23, d39);
	buf (d106, d61);
	not (d107, d8);
	nor (d108, d19, d72);
	nand (d109, d50, d79);
	nand (d110, d26, d78);
	nor (d111, d46, d92);
	nor (d112, d30, d60);
	xor (d113, d55, d70);
	or (d114, d75, d77);
	nor (d115, d77, d87);
	or (d116, d67, d85);
	or (d117, d84, d86);
	nand (d118, d43, d64);
	xor (d119, d27, d96);
	nor (d120, d75, d78);
	and (d121, d44, d74);
	xor (d122, d69, d79);
	xnor (d123, d72, d93);
	nor (d124, d53, d58);
	nor (d125, d57, d90);
	or (d126, d39, d74);
	nor (d127, d52, d74);
	nor (d128, d79, d91);
	nand (d129, d68, d80);
	or (d130, d18, d53);
	or (d131, d28, d43);
	xor (d132, d43, d64);
	not (d133, d94);
	nand (d134, d65, d96);
	and (d135, d30, d82);
	nand (d136, d26, d44);
	xnor (d137, d40, d64);
	xnor (d138, d26, d93);
	nand (d139, d26, d70);
	not (d140, d51);
	nor (d141, d32, d37);
	buf (d142, d60);
	or (d143, d51, d60);
	or (d144, d19, d94);
	and (d145, d28, d74);
	buf (d146, d78);
	and (d147, d56, d84);
	not (d148, d76);
	xnor (d149, d32, d47);
	nand (d150, d63, d91);
	buf (d151, d10);
	not (d152, d55);
	buf (d153, d3);
	buf (d154, d32);
	or (d155, d59, d78);
	or (d156, d22, d53);
	xnor (d157, d50, d53);
	assign f1 = d116;
	assign f2 = d115;
	assign f3 = d121;
	assign f4 = d109;
	assign f5 = d99;
	assign f6 = d132;
	assign f7 = d111;
	assign f8 = d149;
	assign f9 = d123;
	assign f10 = d150;
	assign f11 = d119;
	assign f12 = d141;
endmodule
