module CCGRCG82( x0, x1, x2, x3, f1, f2, f3, f4, f5 );

	input x0, x1, x2, x3;
	output f1, f2, f3, f4, f5;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314, d315, d316, d317, d318, d319, d320, d321, d322;

	not (d1, x2);
	or (d2, x1, x3);
	xor (d3, x0, x2);
	nor (d4, x3);
	nand (d5, x0, x3);
	not (d6, x3);
	not (d7, x0);
	or (d8, x0);
	xnor (d9, x2, x3);
	xnor (d10, x0, x2);
	or (d11, x3);
	and (d12, x0, x2);
	and (d13, x1, x3);
	xnor (d14, x0);
	nor (d15, x2);
	xor (d16, x0);
	xnor (d17, x1, x2);
	xor (d18, x2, x3);
	or (d19, x1, x3);
	not (d20, x1);
	buf (d21, x1);
	xor (d22, x1, x2);
	nor (d23, x2, x3);
	or (d24, x0, x2);
	or (d25, x0, x1);
	nand (d26, x2, x3);
	buf (d27, x2);
	and (d28, x0, x3);
	nand (d29, x1, x2);
	nand (d30, x0);
	xor (d31, d20, d29);
	and (d32, d9, d19);
	xor (d33, d15, d24);
	not (d34, d28);
	nand (d35, d16, d20);
	nor (d36, d20);
	or (d37, d9, d15);
	nor (d38, d9, d28);
	xor (d39, d27, d28);
	xnor (d40, d11, d13);
	buf (d41, d11);
	or (d42, d4, d12);
	nor (d43, d8, d29);
	nor (d44, d43);
	nand (d45, d33, d38);
	xnor (d46, d31, d43);
	buf (d47, d42);
	and (d48, d36, d39);
	or (d49, d31, d33);
	xnor (d50, d40, d42);
	nand (d51, d32, d38);
	nor (d52, d35, d40);
	xor (d53, d34, d36);
	nor (d54, d32);
	nor (d55, d31, d37);
	nand (d56, d35, d40);
	nor (d57, d36, d39);
	nor (d58, d41, d43);
	nor (d59, d33, d43);
	xor (d60, d34, d40);
	and (d61, d31, d32);
	not (d62, d19);
	nand (d63, d34, d35);
	not (d64, d12);
	nor (d65, d33, d34);
	not (d66, d14);
	nand (d67, d36, d43);
	xnor (d68, d34, d43);
	nand (d69, d35, d39);
	and (d70, d35, d41);
	xnor (d71, d36, d39);
	and (d72, d36, d43);
	nor (d73, d39, d43);
	nand (d74, d37, d39);
	and (d75, d32, d38);
	nand (d76, d38);
	buf (d77, d26);
	nor (d78, d34, d38);
	not (d79, d38);
	and (d80, d38, d40);
	or (d81, d33, d35);
	xor (d82, d34, d35);
	not (d83, d27);
	xnor (d84, d36, d37);
	not (d85, d40);
	nor (d86, d38, d43);
	xor (d87, d36, d40);
	xor (d88, d35);
	not (d89, d26);
	nand (d90, d33, d39);
	xnor (d91, d33, d40);
	nand (d92, d34);
	nor (d93, d33, d34);
	buf (d94, d16);
	not (d95, d10);
	and (d96, d41);
	or (d97, d35, d41);
	xnor (d98, d36, d41);
	buf (d99, d20);
	xor (d100, d34, d42);
	xor (d101, d37, d42);
	and (d102, d38, d43);
	and (d103, d35, d37);
	and (d104, d36, d43);
	buf (d105, d9);
	and (d106, d32, d39);
	and (d107, d35, d43);
	or (d108, d36, d40);
	nor (d109, d38, d39);
	nand (d110, d32, d37);
	xor (d111, d34, d40);
	and (d112, d37, d38);
	xnor (d113, d35, d41);
	and (d114, d32);
	and (d115, d33, d38);
	and (d116, d31, d36);
	xor (d117, d39, d43);
	nor (d118, d32, d33);
	buf (d119, d29);
	not (d120, d21);
	xor (d121, d31, d38);
	or (d122, d39);
	xnor (d123, d35, d43);
	or (d124, d32, d39);
	or (d125, d34, d39);
	or (d126, d32, d33);
	buf (d127, d1);
	not (d128, d43);
	not (d129, d39);
	xor (d130, d35, d40);
	nand (d131, d36, d41);
	not (d132, d4);
	nand (d133, d40, d43);
	not (d134, d30);
	buf (d135, d53);
	buf (d136, d133);
	buf (d137, d4);
	and (d138, d46, d75);
	or (d139, d51, d129);
	nor (d140, d47, d128);
	nand (d141, d55, d77);
	xor (d142, d45, d119);
	not (d143, d24);
	nor (d144, d105, d127);
	buf (d145, d57);
	or (d146, d64, d121);
	not (d147, d89);
	buf (d148, d103);
	and (d149, d57, d98);
	xnor (d150, d63, d83);
	or (d151, d90, d130);
	not (d152, d59);
	nor (d153, d93, d122);
	not (d154, d41);
	not (d155, d105);
	xor (d156, d69, d92);
	xnor (d157, d48, d50);
	xor (d158, d85, d126);
	and (d159, d66, d72);
	xor (d160, d76, d85);
	nand (d161, d123, d124);
	nor (d162, d80, d86);
	xor (d163, d105, d134);
	xor (d164, d75, d125);
	xnor (d165, d64, d86);
	xnor (d166, d54, d57);
	xnor (d167, d106, d132);
	xor (d168, d70, d87);
	and (d169, d119, d125);
	nor (d170, d72, d117);
	and (d171, d59, d106);
	nor (d172, d68, d98);
	xnor (d173, d55, d119);
	nand (d174, d46, d92);
	not (d175, d107);
	xor (d176, d70, d90);
	xor (d177, d80, d114);
	xnor (d178, d56, d124);
	and (d179, d58, d128);
	buf (d180, d117);
	xnor (d181, d72, d120);
	and (d182, d53, d75);
	not (d183, d101);
	nand (d184, d105, d128);
	nor (d185, d59, d103);
	xnor (d186, d84, d128);
	nor (d187, d51, d98);
	nand (d188, d65, d89);
	buf (d189, d63);
	nand (d190, d79, d129);
	and (d191, d84, d123);
	and (d192, d79, d104);
	and (d193, d131, d134);
	buf (d194, d94);
	xor (d195, d53, d89);
	xor (d196, d45, d67);
	buf (d197, d116);
	and (d198, d107, d112);
	buf (d199, d56);
	nor (d200, d61, d71);
	not (d201, d130);
	nand (d202, d105);
	nand (d203, d47, d55);
	nand (d204, d70, d96);
	and (d205, d57, d130);
	nor (d206, d75, d104);
	xor (d207, d144, d188);
	nand (d208, d155, d190);
	nor (d209, d158, d195);
	nand (d210, d148, d152);
	xnor (d211, d178, d198);
	not (d212, d48);
	or (d213, d181, d189);
	nand (d214, d144, d181);
	not (d215, d42);
	nand (d216, d135, d161);
	not (d217, d153);
	or (d218, d139, d195);
	buf (d219, d149);
	nand (d220, d157, d162);
	xor (d221, d141, d183);
	not (d222, d167);
	xor (d223, d188, d198);
	nor (d224, d144, d183);
	xnor (d225, d146, d188);
	and (d226, d137, d175);
	buf (d227, d168);
	nor (d228, d175, d201);
	nand (d229, d165, d176);
	xnor (d230, d143, d202);
	xor (d231, d165, d182);
	or (d232, d159, d166);
	nand (d233, d216, d227);
	xnor (d234, d214, d215);
	or (d235, d222, d224);
	xor (d236, d217, d220);
	nor (d237, d211, d229);
	nor (d238, d208, d225);
	or (d239, d207, d208);
	not (d240, d174);
	xor (d241, d221, d226);
	and (d242, d214, d222);
	buf (d243, d71);
	and (d244, d207, d221);
	xnor (d245, d211, d212);
	xnor (d246, d212, d215);
	buf (d247, d62);
	xnor (d248, d211, d215);
	nor (d249, d224, d231);
	nor (d250, d214, d224);
	and (d251, d208, d223);
	not (d252, d126);
	not (d253, d94);
	buf (d254, d151);
	or (d255, d210, d217);
	buf (d256, d221);
	xor (d257, d216, d222);
	xnor (d258, d209, d212);
	xor (d259, d211, d215);
	and (d260, d210, d231);
	buf (d261, d153);
	buf (d262, d145);
	or (d263, d220, d231);
	not (d264, d18);
	nor (d265, d216, d219);
	nand (d266, d220, d229);
	not (d267, d15);
	nand (d268, d218, d230);
	nor (d269, d208, d218);
	or (d270, d218, d220);
	not (d271, d74);
	xor (d272, d207, d226);
	xnor (d273, d218, d226);
	xor (d274, d210, d220);
	buf (d275, d211);
	buf (d276, d51);
	or (d277, d220);
	nand (d278, d207, d224);
	and (d279, d207, d213);
	xnor (d280, d223, d227);
	or (d281, d217, d227);
	xnor (d282, d211, d218);
	xor (d283, d216, d223);
	not (d284, d215);
	buf (d285, d171);
	xor (d286, d211, d213);
	nand (d287, d209, d210);
	and (d288, d208, d232);
	or (d289, d217, d225);
	not (d290, d68);
	buf (d291, d75);
	and (d292, d212, d232);
	and (d293, d217, d218);
	buf (d294, d201);
	nor (d295, d210, d217);
	nand (d296, d224, d226);
	xor (d297, d208, d225);
	and (d298, d211, d227);
	or (d299, d215, d232);
	nand (d300, d215, d226);
	and (d301, d227, d232);
	nand (d302, d219, d224);
	xor (d303, d216, d220);
	nand (d304, d210, d232);
	buf (d305, d2);
	buf (d306, d88);
	or (d307, d208, d210);
	buf (d308, d3);
	buf (d309, d129);
	nand (d310, d211, d228);
	buf (d311, d30);
	buf (d312, d177);
	nor (d313, d211, d219);
	or (d314, d208, d225);
	nand (d315, d211, d225);
	or (d316, d209, d211);
	xor (d317, d209, d219);
	and (d318, d223, d230);
	xor (d319, d213, d217);
	xor (d320, d209, d213);
	not (d321, d232);
	xnor (d322, d215, d218);
	assign f1 = d310;
	assign f2 = d262;
	assign f3 = d237;
	assign f4 = d269;
	assign f5 = d262;
endmodule
