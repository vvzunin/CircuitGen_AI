module CCGRCG180( x0, x1, x2, x3, x4, x5, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16 );

	input x0, x1, x2, x3, x4, x5;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314, d315, d316, d317, d318, d319, d320, d321, d322, d323, d324, d325, d326, d327, d328, d329, d330, d331, d332, d333, d334, d335, d336, d337, d338, d339, d340, d341, d342, d343, d344, d345, d346, d347, d348, d349, d350, d351, d352, d353, d354, d355, d356, d357, d358, d359, d360, d361, d362, d363, d364, d365, d366, d367, d368, d369, d370, d371, d372, d373, d374, d375, d376, d377, d378, d379, d380, d381, d382, d383, d384, d385, d386, d387, d388, d389, d390, d391, d392, d393, d394, d395, d396, d397, d398, d399, d400, d401, d402, d403, d404, d405, d406, d407, d408, d409, d410, d411, d412, d413, d414, d415, d416, d417, d418, d419, d420, d421, d422, d423, d424, d425, d426, d427, d428, d429, d430, d431, d432, d433, d434, d435, d436, d437, d438, d439, d440, d441, d442, d443, d444, d445, d446, d447, d448, d449, d450, d451, d452, d453, d454, d455, d456, d457, d458, d459, d460, d461, d462, d463, d464, d465, d466, d467, d468, d469, d470, d471, d472, d473, d474, d475, d476, d477, d478, d479, d480, d481, d482, d483, d484, d485, d486, d487, d488, d489, d490, d491, d492, d493, d494, d495, d496, d497, d498, d499, d500, d501, d502, d503, d504, d505, d506, d507, d508, d509, d510, d511, d512, d513, d514, d515, d516, d517, d518, d519, d520, d521, d522, d523, d524, d525, d526, d527, d528, d529, d530, d531, d532, d533, d534, d535, d536, d537, d538, d539, d540, d541, d542, d543, d544, d545, d546, d547, d548, d549, d550, d551, d552, d553;

	nand (d1, x1, x3);
	not (d2, x1);
	or (d3, x1, x5);
	xor (d4, x1, x5);
	xnor (d5, x2, x5);
	nor (d6, x3);
	xor (d7, x1, x3);
	xnor (d8, x0, x3);
	xnor (d9, x3);
	and (d10, x1, x5);
	nand (d11, x1, x5);
	nand (d12, x2, x3);
	or (d13, x0, x5);
	or (d14, x2, x3);
	buf (d15, x0);
	xnor (d16, x1, x3);
	xnor (d17, x1, x5);
	buf (d18, x5);
	and (d19, x0, x2);
	and (d20, x0);
	nand (d21, d4, d12);
	buf (d22, d19);
	xnor (d23, d2, d14);
	buf (d24, d2);
	buf (d25, d1);
	or (d26, d1, d16);
	nand (d27, d6, d7);
	nand (d28, d2, d16);
	buf (d29, d3);
	or (d30, d8, d20);
	or (d31, d4, d18);
	nand (d32, d14, d20);
	xnor (d33, d19, d20);
	xor (d34, d9);
	xor (d35, d12, d19);
	nor (d36, d10, d11);
	not (d37, d18);
	and (d38, d6, d17);
	nor (d39, d8, d16);
	nor (d40, d3, d9);
	or (d41, d5, d6);
	and (d42, d8, d12);
	nor (d43, d2, d13);
	or (d44, d7, d18);
	buf (d45, x2);
	and (d46, d6, d10);
	xnor (d47, d6, d7);
	nor (d48, d3, d16);
	and (d49, d6, d16);
	or (d50, d1, d9);
	xnor (d51, d8, d11);
	nor (d52, d15, d19);
	xnor (d53, d5, d15);
	nand (d54, d14, d15);
	xnor (d55, d8, d11);
	xnor (d56, d5, d6);
	or (d57, d7, d17);
	and (d58, d2, d3);
	nor (d59, d14, d19);
	xor (d60, d10, d15);
	nor (d61, d4, d19);
	xor (d62, d11, d17);
	nor (d63, d18, d19);
	or (d64, d4, d10);
	and (d65, d10, d17);
	nand (d66, d6, d11);
	or (d67, d1, d5);
	or (d68, d1, d9);
	nand (d69, d10, d11);
	xor (d70, d13);
	buf (d71, d13);
	xnor (d72, d18, d20);
	xnor (d73, d15, d19);
	nor (d74, d14, d18);
	buf (d75, d11);
	not (d76, d7);
	xnor (d77, d2, d10);
	xnor (d78, d11, d16);
	nor (d79, d4, d6);
	nor (d80, d5, d16);
	and (d81, d4, d14);
	xor (d82, d11, d18);
	not (d83, d8);
	not (d84, d11);
	and (d85, d8);
	nor (d86, d8, d17);
	buf (d87, d16);
	or (d88, d3, d19);
	xor (d89, d10, d17);
	not (d90, d1);
	xor (d91, d6, d18);
	and (d92, d2, d10);
	xor (d93, d4, d7);
	xnor (d94, d5, d16);
	xor (d95, d1, d5);
	buf (d96, d7);
	or (d97, d5, d11);
	buf (d98, d15);
	xnor (d99, d8, d16);
	xnor (d100, d73, d79);
	buf (d101, d58);
	nor (d102, d22, d62);
	nand (d103, d65, d68);
	xor (d104, d34, d46);
	xnor (d105, d50, d65);
	not (d106, d9);
	not (d107, d78);
	xor (d108, d42, d45);
	xor (d109, d65, d82);
	buf (d110, d81);
	buf (d111, d23);
	or (d112, d56, d82);
	xor (d113, d23, d81);
	xnor (d114, d47, d55);
	buf (d115, d78);
	nand (d116, d50, d65);
	and (d117, d29, d52);
	and (d118, d22, d99);
	or (d119, d56, d58);
	and (d120, d75, d90);
	not (d121, d13);
	not (d122, d75);
	and (d123, d53, d89);
	not (d124, d83);
	not (d125, d22);
	xor (d126, d25, d92);
	nand (d127, d31, d96);
	xnor (d128, d68, d83);
	xnor (d129, d83, d93);
	xnor (d130, d23, d80);
	xnor (d131, d35, d71);
	nand (d132, d32, d84);
	or (d133, d82);
	xor (d134, d118, d130);
	buf (d135, d105);
	xnor (d136, d104, d133);
	and (d137, d112, d120);
	or (d138, d116, d120);
	nand (d139, d100, d112);
	xnor (d140, d102, d128);
	xor (d141, d104, d116);
	or (d142, d125, d133);
	nand (d143, d105, d116);
	nor (d144, d128, d131);
	or (d145, d107, d121);
	not (d146, d30);
	xnor (d147, d110, d112);
	not (d148, d39);
	nor (d149, d104, d111);
	nand (d150, d109, d119);
	nor (d151, d128, d129);
	nand (d152, d106, d125);
	xnor (d153, d120, d122);
	buf (d154, d28);
	nand (d155, d104, d126);
	buf (d156, d91);
	xor (d157, d123, d124);
	and (d158, d111, d133);
	buf (d159, d10);
	xnor (d160, d119, d123);
	and (d161, d113, d122);
	nor (d162, d114, d122);
	nand (d163, d105, d131);
	nand (d164, d130, d132);
	or (d165, d101, d120);
	or (d166, d107, d120);
	buf (d167, d60);
	xnor (d168, d105, d107);
	xor (d169, d111, d112);
	xnor (d170, d105, d109);
	and (d171, d101, d122);
	nand (d172, d107, d110);
	and (d173, d101, d113);
	xnor (d174, d104, d127);
	xnor (d175, d112, d133);
	or (d176, d102, d115);
	not (d177, d123);
	nor (d178, d116, d133);
	xor (d179, d108, d118);
	or (d180, d114, d115);
	or (d181, d100, d128);
	buf (d182, d68);
	buf (d183, d109);
	xnor (d184, d102, d117);
	nor (d185, d103, d115);
	nor (d186, d104, d118);
	and (d187, d105, d112);
	nor (d188, d103, d122);
	xnor (d189, d104, d111);
	nand (d190, d116, d126);
	xor (d191, d112, d122);
	not (d192, d129);
	buf (d193, d55);
	xor (d194, d104, d121);
	nand (d195, d114, d126);
	nand (d196, d101, d106);
	nor (d197, d106, d113);
	xnor (d198, d106, d127);
	nand (d199, d102, d115);
	not (d200, d122);
	buf (d201, d64);
	nor (d202, d127, d132);
	and (d203, d119, d123);
	nand (d204, d100, d129);
	xor (d205, d115, d132);
	nand (d206, d106, d124);
	xor (d207, d122, d125);
	xnor (d208, d105, d132);
	and (d209, d110, d122);
	xor (d210, d115, d119);
	xor (d211, d114, d129);
	not (d212, d126);
	buf (d213, d79);
	xor (d214, d119, d127);
	xor (d215, d111, d113);
	nor (d216, d100, d114);
	xor (d217, d128, d131);
	xnor (d218, d102, d118);
	and (d219, d119, d127);
	and (d220, d100, d107);
	nand (d221, d106, d108);
	and (d222, d101, d120);
	and (d223, d102, d113);
	xnor (d224, d104, d123);
	and (d225, d179, d191);
	buf (d226, d150);
	xor (d227, d187, d206);
	and (d228, d134, d167);
	buf (d229, d219);
	xnor (d230, d174, d180);
	nor (d231, d188, d192);
	nor (d232, d135, d175);
	not (d233, d216);
	xnor (d234, d200, d212);
	xor (d235, d150, d203);
	or (d236, d179, d209);
	not (d237, d91);
	nor (d238, d170, d174);
	xor (d239, d171, d181);
	not (d240, d193);
	nand (d241, d135, d177);
	nor (d242, d143, d158);
	xor (d243, d188, d224);
	xor (d244, d137, d200);
	or (d245, d137, d156);
	xnor (d246, d167, d213);
	nor (d247, d184, d205);
	and (d248, d135, d190);
	nand (d249, d145, d206);
	not (d250, d155);
	not (d251, d85);
	and (d252, d154, d208);
	not (d253, d69);
	buf (d254, d171);
	not (d255, d177);
	and (d256, d162, d200);
	xor (d257, d183, d213);
	xor (d258, d173, d213);
	buf (d259, d88);
	nor (d260, d147, d181);
	and (d261, d208, d217);
	nor (d262, d145, d183);
	xnor (d263, d152, d195);
	and (d264, d167, d220);
	or (d265, d193, d198);
	buf (d266, d152);
	buf (d267, d114);
	or (d268, d141, d206);
	nor (d269, d136, d138);
	not (d270, d32);
	or (d271, d149, d153);
	or (d272, d146, d214);
	or (d273, d154, d171);
	xor (d274, d138, d187);
	or (d275, d162, d209);
	or (d276, d144, d153);
	nand (d277, d141, d162);
	and (d278, d140, d164);
	nand (d279, d141, d211);
	and (d280, d163, d196);
	or (d281, d183, d189);
	or (d282, d142, d178);
	xor (d283, d149, d214);
	xor (d284, d153, d203);
	buf (d285, d143);
	nand (d286, d151, d167);
	or (d287, d197, d222);
	nand (d288, d161, d185);
	buf (d289, d83);
	nand (d290, d197, d208);
	xnor (d291, d165, d206);
	buf (d292, d5);
	and (d293, d144, d187);
	nand (d294, d156, d171);
	buf (d295, d214);
	buf (d296, d26);
	or (d297, d144, d203);
	buf (d298, d170);
	buf (d299, d97);
	nand (d300, d172, d200);
	not (d301, d55);
	and (d302, d149, d224);
	nor (d303, d142, d208);
	or (d304, d192, d216);
	or (d305, d152);
	nand (d306, d283, d299);
	nand (d307, d247, d269);
	not (d308, d79);
	nand (d309, d289, d290);
	nand (d310, d225, d249);
	or (d311, d239, d263);
	or (d312, d227, d260);
	not (d313, d218);
	or (d314, d251, d252);
	or (d315, d278, d297);
	nor (d316, d241, d244);
	xor (d317, d258, d284);
	nand (d318, d230, d261);
	xnor (d319, d250, d258);
	not (d320, d66);
	and (d321, d271, d290);
	and (d322, d264, d303);
	nand (d323, d255, d256);
	xor (d324, d251, d262);
	and (d325, d249, d295);
	xor (d326, d244, d300);
	and (d327, d277, d300);
	buf (d328, d217);
	not (d329, d130);
	and (d330, d238, d264);
	nand (d331, d248, d264);
	or (d332, d231, d294);
	nand (d333, d262, d300);
	nor (d334, d234, d238);
	and (d335, d265, d300);
	not (d336, d298);
	xor (d337, d286, d296);
	and (d338, d225, d260);
	not (d339, d180);
	nand (d340, d242, d249);
	buf (d341, d45);
	xor (d342, d250, d269);
	not (d343, d285);
	xor (d344, d248, d299);
	nand (d345, d255, d300);
	or (d346, d244, d304);
	or (d347, d232, d285);
	xnor (d348, d256, d280);
	or (d349, d228, d289);
	xor (d350, d259, d286);
	xor (d351, d286, d295);
	xor (d352, d236, d284);
	or (d353, d248, d259);
	buf (d354, d141);
	nor (d355, d273, d283);
	nand (d356, d259, d275);
	xnor (d357, d229, d246);
	xor (d358, d244, d259);
	nor (d359, d272, d286);
	nor (d360, d227, d242);
	xor (d361, d245, d287);
	xnor (d362, d228, d250);
	xor (d363, d244, d298);
	and (d364, d259, d295);
	nand (d365, d234, d297);
	xnor (d366, d325, d362);
	or (d367, d316, d353);
	or (d368, d344, d351);
	xor (d369, d324, d356);
	or (d370, d348, d360);
	xnor (d371, d341, d353);
	buf (d372, d304);
	xnor (d373, d307, d364);
	nor (d374, d334, d340);
	xor (d375, d316, d345);
	xnor (d376, d317, d353);
	nor (d377, d330);
	not (d378, d319);
	xnor (d379, d306, d348);
	xor (d380, d309, d342);
	buf (d381, d75);
	or (d382, d326, d341);
	xnor (d383, d342, d365);
	not (d384, d206);
	buf (d385, d360);
	or (d386, d354, d361);
	xor (d387, d333, d347);
	or (d388, d339, d359);
	not (d389, d286);
	or (d390, d308, d355);
	nand (d391, d347, d349);
	not (d392, d35);
	xor (d393, d356, d362);
	not (d394, d301);
	nor (d395, d353, d354);
	buf (d396, d317);
	buf (d397, d359);
	xor (d398, d375, d395);
	xnor (d399, d389, d394);
	and (d400, d377, d393);
	or (d401, d366, d373);
	nand (d402, d380, d381);
	not (d403, d333);
	xor (d404, d388, d392);
	buf (d405, d338);
	xor (d406, d367, d383);
	nand (d407, d387, d389);
	nand (d408, d370, d391);
	buf (d409, d309);
	not (d410, d304);
	or (d411, d377, d389);
	nor (d412, d382, d391);
	or (d413, d376, d382);
	not (d414, d339);
	nor (d415, d371, d375);
	xnor (d416, d371, d393);
	xor (d417, d377, d382);
	nand (d418, d388, d394);
	and (d419, d371, d395);
	nand (d420, d378, d386);
	xor (d421, d377, d390);
	buf (d422, d12);
	or (d423, d390, d394);
	nor (d424, d377, d380);
	xnor (d425, d377, d379);
	nor (d426, d384, d386);
	nand (d427, d379, d391);
	nand (d428, d379, d382);
	and (d429, d380, d388);
	and (d430, d386, d390);
	buf (d431, d140);
	not (d432, d237);
	not (d433, d113);
	buf (d434, d267);
	xor (d435, d391, d392);
	and (d436, d381, d383);
	not (d437, d313);
	xnor (d438, d378, d384);
	buf (d439, d221);
	or (d440, d390, d391);
	xnor (d441, d387, d388);
	and (d442, d385, d387);
	xnor (d443, d367, d372);
	nor (d444, d374, d385);
	xnor (d445, d373, d392);
	nand (d446, d371, d373);
	nor (d447, d388, d391);
	or (d448, d370, d394);
	xor (d449, d380, d381);
	nor (d450, d366, d376);
	or (d451, d374, d378);
	not (d452, d179);
	xor (d453, d374, d383);
	nand (d454, d382, d391);
	nor (d455, d390, d393);
	or (d456, d368, d374);
	nor (d457, d380, d395);
	xnor (d458, d374, d381);
	and (d459, d387, d390);
	xor (d460, d366, d380);
	xor (d461, d389, d395);
	not (d462, d198);
	not (d463, d280);
	or (d464, d381, d387);
	xor (d465, d376, d384);
	xor (d466, d381, d382);
	xor (d467, d381, d391);
	buf (d468, d40);
	or (d469, d369, d388);
	or (d470, d378, d386);
	nor (d471, d389, d390);
	or (d472, d433, d451);
	nor (d473, d461, d471);
	nand (d474, d413, d467);
	nor (d475, d446, d457);
	nand (d476, d424, d457);
	nand (d477, d403, d454);
	and (d478, d435, d462);
	nand (d479, d446, d457);
	not (d480, d471);
	and (d481, d420, d441);
	nor (d482, d447, d457);
	xnor (d483, d406, d427);
	xor (d484, d404, d439);
	xnor (d485, d398, d471);
	buf (d486, d257);
	and (d487, d397, d465);
	nor (d488, d419, d461);
	nand (d489, d442, d466);
	or (d490, d397, d430);
	nor (d491, d427, d469);
	or (d492, d430, d438);
	not (d493, d252);
	buf (d494, d436);
	xor (d495, d442, d460);
	xor (d496, d436, d442);
	xor (d497, d450, d463);
	xor (d498, d400, d411);
	not (d499, d306);
	and (d500, d436, d464);
	nor (d501, d425, d469);
	nor (d502, d402, d405);
	xnor (d503, d406, d429);
	and (d504, d396, d452);
	not (d505, d139);
	xor (d506, d397, d420);
	buf (d507, d256);
	not (d508, d184);
	and (d509, d421, d427);
	not (d510, d53);
	xor (d511, d457, d461);
	xor (d512, d435, d455);
	xor (d513, d396, d449);
	nor (d514, d401, d439);
	or (d515, d422, d466);
	nand (d516, d409, d419);
	xor (d517, d444, d465);
	nor (d518, d445, d448);
	not (d519, d341);
	not (d520, d136);
	and (d521, d435, d458);
	xor (d522, d453, d462);
	and (d523, d453, d465);
	nand (d524, d408, d412);
	nand (d525, d441, d456);
	or (d526, d400, d409);
	buf (d527, d85);
	buf (d528, d76);
	and (d529, d433, d469);
	nor (d530, d418, d436);
	xnor (d531, d398, d427);
	xor (d532, d397, d459);
	not (d533, d14);
	nor (d534, d397, d437);
	and (d535, d421, d469);
	xor (d536, d427, d449);
	not (d537, d365);
	and (d538, d431, d456);
	buf (d539, d397);
	xnor (d540, d423, d453);
	buf (d541, d207);
	and (d542, d424, d455);
	xnor (d543, d412, d445);
	xnor (d544, d428, d464);
	buf (d545, d192);
	xnor (d546, d443, d459);
	xor (d547, d422, d435);
	xnor (d548, d462, d470);
	nand (d549, d420, d469);
	or (d550, d453, d455);
	and (d551, d438, d456);
	xnor (d552, d420, d464);
	xnor (d553, d432, d448);
	assign f1 = d506;
	assign f2 = d515;
	assign f3 = d515;
	assign f4 = d493;
	assign f5 = d507;
	assign f6 = d520;
	assign f7 = d527;
	assign f8 = d472;
	assign f9 = d537;
	assign f10 = d521;
	assign f11 = d521;
	assign f12 = d515;
	assign f13 = d492;
	assign f14 = d496;
	assign f15 = d552;
	assign f16 = d519;
endmodule
