module CCGRCG6( x0, x1, f1, f2, f3, f4, f5 );

	input x0, x1;
	output f1, f2, f3, f4, f5;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62;

	nor (d1, x0, x1);
	or (d2, x0, x1);
	and (d3, x0);
	nor (d4, x0, x1);
	not (d5, x1);
	or (d6, d1);
	xor (d7, d2, d5);
	buf (d8, x0);
	or (d9, d3, d4);
	or (d10, d2, d4);
	not (d11, x0);
	or (d12, d4, d5);
	buf (d13, x1);
	nor (d14, d2, d5);
	not (d15, d3);
	xor (d16, d1, d5);
	nand (d17, d4, d5);
	nor (d18, d5);
	xor (d19, d1, d2);
	and (d20, d2, d4);
	buf (d21, d5);
	nor (d22, d1, d4);
	xor (d23, d2, d3);
	xor (d24, d1, d4);
	xor (d25, d2, d5);
	or (d26, d3, d5);
	buf (d27, d3);
	or (d28, d2, d5);
	nand (d29, d1, d3);
	nand (d30, d1, d3);
	xor (d31, d5);
	not (d32, d1);
	nand (d33, d3, d5);
	nand (d34, d2, d3);
	not (d35, d5);
	and (d36, d1, d5);
	nor (d37, d4, d5);
	xor (d38, d1, d3);
	or (d39, d4);
	nand (d40, d3, d4);
	xnor (d41, d2, d4);
	nand (d42, d4);
	and (d43, d3);
	or (d44, d3);
	xor (d45, d4, d5);
	xnor (d46, d4, d5);
	buf (d47, d1);
	nand (d48, d3);
	xnor (d49, d3, d4);
	xor (d50, d2);
	or (d51, d2, d3);
	and (d52, d2, d3);
	nand (d53, d4, d5);
	and (d54, d2, d5);
	not (d55, d2);
	and (d56, d4);
	nand (d57, d5);
	nand (d58, d1, d2);
	nand (d59, d2, d4);
	xor (d60, d2, d4);
	xnor (d61, d2);
	or (d62, d1, d4);
	assign f1 = d37;
	assign f2 = d45;
	assign f3 = d13;
	assign f4 = d27;
	assign f5 = d13;
endmodule
