module CCGRCG185( x0, x1, x2, x3, x4, x5, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17, f18 );

	input x0, x1, x2, x3, x4, x5;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17, f18;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40;

	and (d1, x2, x5);
	or (d2, x1, x4);
	xor (d3, x1, x3);
	and (d4, x0, x2);
	buf (d5, x2);
	nand (d6, x0, x5);
	not (d7, x2);
	and (d8, x5);
	xnor (d9, x3, x5);
	xnor (d10, x1, x3);
	not (d11, x4);
	nand (d12, x1, x5);
	xnor (d13, x0, x4);
	nor (d14, x3, x5);
	nor (d15, x0, x1);
	xor (d16, x3, x4);
	xnor (d17, x1);
	xor (d18, x3, x5);
	and (d19, x2, x3);
	not (d20, x3);
	nor (d21, x1, x5);
	nor (d22, x5);
	not (d23, x1);
	xnor (d24, x2, x3);
	or (d25, x2, x4);
	xnor (d26, x1, x4);
	and (d27, x4);
	buf (d28, x5);
	or (d29, x4);
	and (d30, x4, x5);
	nor (d31, x4, x5);
	nand (d32, x1, x5);
	or (d33, x2, x5);
	nor (d34, x1, x2);
	and (d35, x0, x4);
	or (d36, x0, x5);
	xnor (d37, x1, x5);
	and (d38, x3, x4);
	nor (d39, x3);
	xnor (d40, x0, x1);
	assign f1 = d10;
	assign f2 = d7;
	assign f3 = d35;
	assign f4 = d4;
	assign f5 = d32;
	assign f6 = d28;
	assign f7 = d1;
	assign f8 = d28;
	assign f9 = d24;
	assign f10 = d2;
	assign f11 = d19;
	assign f12 = d40;
	assign f13 = d39;
	assign f14 = d6;
	assign f15 = d27;
	assign f16 = d20;
	assign f17 = d17;
	assign f18 = d7;
endmodule
