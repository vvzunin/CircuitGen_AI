module CCGRCG69( x0, x1, x2, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17 );

	input x0, x1, x2;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146;

	xnor (d1, x0, x1);
	and (d2, x1, x2);
	or (d3, x1, x2);
	nor (d4, x0, x2);
	nor (d5, x0, x1);
	nand (d6, x1, x2);
	buf (d7, x0);
	and (d8, x0, x2);
	not (d9, x1);
	or (d10, x0, x2);
	and (d11, x0);
	xnor (d12, x1, x2);
	or (d13, x0, x1);
	not (d14, x2);
	or (d15, x0, x1);
	xnor (d16, x0, x1);
	nand (d17, x0, x1);
	nor (d18, x1, x2);
	xor (d19, x0, x1);
	or (d20, x0, x2);
	xor (d21, x0);
	nand (d22, x2);
	xor (d23, x0, x2);
	and (d24, x2);
	and (d25, x0, x2);
	buf (d26, x1);
	nand (d27, x1, x2);
	buf (d28, x2);
	and (d29, x1);
	not (d30, x0);
	xor (d31, x0, x1);
	xnor (d32, x1);
	xnor (d33, x0, x2);
	nor (d34, x1);
	xnor (d35, x1, x2);
	nor (d36, x0);
	nor (d37, x0, x2);
	xor (d38, x1, x2);
	xnor (d39, x0, x2);
	xnor (d40, d32, d38);
	buf (d41, d15);
	not (d42, d25);
	or (d43, d2, d15);
	or (d44, d7, d32);
	not (d45, d22);
	xnor (d46, d10, d11);
	buf (d47, d2);
	not (d48, d19);
	nor (d49, d7, d16);
	not (d50, d33);
	nor (d51, d26, d36);
	nand (d52, d30, d33);
	nor (d53, d8, d29);
	nand (d54, d18, d34);
	xor (d55, d19, d24);
	xnor (d56, d15, d21);
	nand (d57, d3, d24);
	xnor (d58, d42, d57);
	xor (d59, d51, d56);
	not (d60, d47);
	xor (d61, d46, d47);
	xnor (d62, d40, d57);
	xnor (d63, d49, d50);
	xnor (d64, d40, d43);
	xnor (d65, d41, d44);
	or (d66, d41, d44);
	nand (d67, d46, d47);
	not (d68, d14);
	nor (d69, d41, d53);
	buf (d70, d5);
	nand (d71, d42, d56);
	nor (d72, d53, d54);
	buf (d73, d51);
	nor (d74, d40, d50);
	or (d75, d43, d57);
	and (d76, d41, d42);
	and (d77, d49, d50);
	buf (d78, d23);
	xnor (d79, d42, d48);
	nand (d80, d41, d46);
	and (d81, d47, d51);
	nand (d82, d45, d56);
	xor (d83, d44, d55);
	xor (d84, d48, d55);
	nand (d85, d48, d56);
	or (d86, d44, d55);
	not (d87, d53);
	buf (d88, d44);
	xnor (d89, d43, d57);
	nor (d90, d44, d57);
	buf (d91, d37);
	buf (d92, d31);
	not (d93, d27);
	nand (d94, d44, d47);
	buf (d95, d43);
	buf (d96, d22);
	nor (d97, d51, d56);
	not (d98, d15);
	not (d99, d24);
	xor (d100, d47, d49);
	xor (d101, d42, d56);
	or (d102, d41, d54);
	or (d103, d53);
	xor (d104, d51, d57);
	nor (d105, d50, d51);
	and (d106, d51, d57);
	or (d107, d42, d53);
	xor (d108, d55, d56);
	xnor (d109, d40, d41);
	and (d110, d55, d56);
	nor (d111, d42, d51);
	nand (d112, d42, d49);
	nand (d113, d55);
	nor (d114, d47, d56);
	xnor (d115, d48, d55);
	or (d116, d45, d53);
	and (d117, d41);
	xnor (d118, d42, d44);
	nand (d119, d54, d57);
	xnor (d120, d42, d54);
	or (d121, d43, d53);
	buf (d122, d49);
	or (d123, d44, d54);
	or (d124, d50, d55);
	xnor (d125, d52, d57);
	nor (d126, d42, d55);
	nand (d127, d42, d53);
	xor (d128, d58, d120);
	buf (d129, d86);
	nor (d130, d120);
	nor (d131, d102, d127);
	xor (d132, d64, d91);
	xnor (d133, d59, d69);
	or (d134, d62, d93);
	nand (d135, d91, d126);
	buf (d136, d101);
	or (d137, d86, d117);
	nand (d138, d87, d115);
	xnor (d139, d67, d75);
	nand (d140, d60, d126);
	nor (d141, d61, d62);
	buf (d142, d88);
	xnor (d143, d71, d107);
	xor (d144, d63, d66);
	nor (d145, d67, d74);
	buf (d146, d82);
	assign f1 = d128;
	assign f2 = d143;
	assign f3 = d137;
	assign f4 = d133;
	assign f5 = d138;
	assign f6 = d143;
	assign f7 = d136;
	assign f8 = d139;
	assign f9 = d145;
	assign f10 = d142;
	assign f11 = d142;
	assign f12 = d135;
	assign f13 = d146;
	assign f14 = d145;
	assign f15 = d137;
	assign f16 = d132;
	assign f17 = d133;
endmodule
