module CCGRCG41( x0, x1, x2, x3, f1 );

	input x0, x1, x2, x3;
	output f1;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143;

	xnor (d1, x1, x3);
	buf (d2, x3);
	and (d3, x1);
	or (d4, x0);
	nor (d5, x0, x1);
	not (d6, x1);
	nor (d7, x1, x3);
	nand (d8, x0, x3);
	and (d9, x2, x3);
	buf (d10, x1);
	and (d11, x0);
	xnor (d12, x2);
	xor (d13, x1, x3);
	nand (d14, x0);
	nand (d15, x3);
	or (d16, x0, x3);
	xor (d17, x0, x1);
	not (d18, x3);
	xnor (d19, x1, x3);
	not (d20, x2);
	nand (d21, x0, x1);
	or (d22, x3);
	nor (d23, x2, x3);
	xor (d24, x1, x2);
	xnor (d25, x1, x2);
	nor (d26, x0, x3);
	buf (d27, x0);
	xnor (d28, x0);
	or (d29, x1, x2);
	nor (d30, x1);
	nand (d31, x0, x2);
	or (d32, x0, x3);
	or (d33, x1, x3);
	xnor (d34, x3);
	or (d35, x0, x2);
	and (d36, x0, x1);
	xnor (d37, d23, d35);
	and (d38, d11, d15);
	xnor (d39, d5, d22);
	xor (d40, d6, d31);
	buf (d41, d5);
	buf (d42, d23);
	nor (d43, d3, d35);
	or (d44, d4, d30);
	buf (d45, x2);
	and (d46, d1, d24);
	buf (d47, d2);
	buf (d48, d13);
	xor (d49, d35);
	or (d50, d21, d36);
	or (d51, d29, d35);
	xnor (d52, d9, d35);
	and (d53, d10, d31);
	xor (d54, d4, d18);
	nor (d55, d30);
	not (d56, d26);
	buf (d57, d31);
	or (d58, d12, d13);
	nand (d59, d13, d17);
	buf (d60, d28);
	xor (d61, d15, d36);
	buf (d62, d9);
	nand (d63, d2, d25);
	and (d64, d19, d20);
	xnor (d65, d18, d27);
	nor (d66, d10, d19);
	xnor (d67, d6, d8);
	and (d68, d1, d10);
	nand (d69, d7, d17);
	and (d70, d32, d33);
	not (d71, d34);
	xnor (d72, d13, d35);
	or (d73, d7, d11);
	and (d74, d4, d11);
	and (d75, d19, d21);
	nand (d76, d13, d26);
	not (d77, d29);
	nor (d78, d8, d36);
	buf (d79, d26);
	nor (d80, d6, d20);
	or (d81, d17, d28);
	and (d82, d2, d24);
	not (d83, d4);
	xnor (d84, d12, d22);
	nor (d85, d6, d16);
	and (d86, d17, d33);
	xor (d87, d4, d30);
	nor (d88, d26, d27);
	or (d89, d2, d31);
	buf (d90, d24);
	nand (d91, d7, d8);
	xnor (d92, d16, d17);
	xor (d93, d14, d23);
	and (d94, d7, d16);
	and (d95, d24, d34);
	not (d96, d25);
	buf (d97, d14);
	xnor (d98, d6, d17);
	nor (d99, d10, d14);
	not (d100, d12);
	and (d101, d8, d27);
	nand (d102, d26, d30);
	xnor (d103, d21, d24);
	buf (d104, d65);
	or (d105, d38, d98);
	not (d106, d14);
	buf (d107, d95);
	nand (d108, d48, d95);
	or (d109, d54, d77);
	xnor (d110, d39, d41);
	or (d111, d66, d81);
	or (d112, d42, d43);
	not (d113, d54);
	or (d114, d37, d97);
	xor (d115, d46, d53);
	nor (d116, d46, d49);
	nand (d117, d40, d97);
	not (d118, d17);
	not (d119, d52);
	not (d120, d68);
	and (d121, d47, d77);
	buf (d122, d8);
	and (d123, d69, d96);
	and (d124, d43, d60);
	xnor (d125, d85);
	nor (d126, d44, d52);
	nor (d127, d56, d102);
	or (d128, d96, d100);
	nand (d129, d43, d103);
	nand (d130, d68, d103);
	xnor (d131, d88, d99);
	not (d132, d42);
	xor (d133, d47, d63);
	buf (d134, d84);
	or (d135, d57, d80);
	xnor (d136, d61, d69);
	not (d137, d40);
	nand (d138, d39, d44);
	not (d139, d90);
	nor (d140, d54, d60);
	or (d141, d51, d69);
	and (d142, d39, d81);
	or (d143, d47, d55);
	assign f1 = d133;
endmodule
