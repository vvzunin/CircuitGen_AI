// Benchmark "CCGRCG128" written by ABC on Tue Feb 13 20:51:59 2024

module CCGRCG128 ( 
    x0, x1, x2, x3, x4,
    f1, f2, f3, f4, f5, f6, f7, f8, f9  );
  input  x0, x1, x2, x3, x4;
  output f1, f2, f3, f4, f5, f6, f7, f8, f9;
  wire new_n16_, new_n17_, new_n19_, new_n20_, new_n21_, new_n22_, new_n23_,
    new_n24_, new_n25_, new_n26_, new_n27_, new_n28_, new_n29_, new_n30_,
    new_n31_, new_n32_, new_n33_, new_n34_, new_n35_, new_n36_, new_n37_,
    new_n38_, new_n39_, new_n40_, new_n41_, new_n42_, new_n43_, new_n44_,
    new_n45_, new_n46_, new_n47_, new_n48_, new_n50_, new_n51_, new_n52_,
    new_n53_, new_n54_, new_n55_, new_n56_, new_n57_, new_n58_, new_n59_,
    new_n60_, new_n62_, new_n63_, new_n64_, new_n65_, new_n66_, new_n67_,
    new_n68_, new_n69_, new_n70_, new_n71_, new_n72_, new_n75_;
  assign new_n16_ = ~x0;
  assign new_n17_ = ~x2;
  assign f8 = ~new_n16_ & ~new_n17_;
  assign new_n19_ = ~x2 & ~x4;
  assign new_n20_ = ~x0 | ~x2;
  assign new_n21_ = new_n20_ ^ new_n19_;
  assign new_n22_ = x3 & x4;
  assign new_n23_ = x1 ^ ~x2;
  assign new_n24_ = ~x1;
  assign new_n25_ = ~x3;
  assign new_n26_ = ~new_n25_ | ~new_n16_ | ~new_n24_;
  assign new_n27_ = ~x1 | (~x0 & ~x3);
  assign new_n28_ = ~new_n26_ | ~new_n27_;
  assign new_n29_ = ~new_n22_ | ~new_n28_ | ~new_n23_;
  assign new_n30_ = ~new_n24_ | ~x2;
  assign new_n31_ = x2 | ~x1;
  assign new_n32_ = ~new_n22_ | ~new_n30_ | ~new_n31_;
  assign new_n33_ = ~new_n27_ | ~new_n32_ | ~new_n26_;
  assign new_n34_ = ~new_n29_ | ~new_n33_;
  assign new_n35_ = ~new_n21_ & ~new_n34_;
  assign new_n36_ = ~new_n35_;
  assign new_n37_ = ~new_n16_ | ~x2;
  assign new_n38_ = x2 | ~x0;
  assign new_n39_ = ~new_n24_ & ~new_n25_;
  assign new_n40_ = ~new_n39_ & (~new_n37_ | ~new_n38_ | ~new_n25_);
  assign new_n41_ = ~x0 & x1;
  assign new_n42_ = new_n19_ | (~new_n17_ & ~new_n41_);
  assign new_n43_ = new_n42_ ? (new_n40_ ^ new_n34_) : (~new_n40_ ^ new_n34_);
  assign new_n44_ = ~x3 | ~x2 | ~new_n24_ | ~x0;
  assign new_n45_ = new_n44_ ^ ~new_n34_;
  assign new_n46_ = ~new_n45_ | ~new_n43_ | ~new_n36_;
  assign new_n47_ = ~new_n46_ | ~f8;
  assign new_n48_ = ~new_n45_ | ~new_n36_ | ~new_n43_ | ~new_n20_;
  assign f2 = ~new_n47_ | ~new_n48_;
  assign new_n50_ = ~new_n43_ | ~new_n36_;
  assign new_n51_ = ~x4;
  assign new_n52_ = ~x2 & ~x3;
  assign new_n53_ = ~new_n20_ | ~new_n44_ | (~new_n51_ & ~new_n52_);
  assign new_n54_ = ~new_n40_;
  assign new_n55_ = ~new_n34_ | ~new_n54_;
  assign new_n56_ = ~new_n40_ | ~new_n29_ | ~new_n33_;
  assign new_n57_ = ~new_n56_ | new_n42_ | ~new_n55_;
  assign new_n58_ = ~new_n55_ | ~new_n56_;
  assign new_n59_ = ~new_n58_ | ~new_n42_;
  assign new_n60_ = ~new_n57_ | ~new_n59_ | ~new_n35_;
  assign f3 = ~new_n53_ & (~new_n50_ | ~new_n60_);
  assign new_n62_ = ~x1 & ~new_n16_;
  assign new_n63_ = ~new_n41_ & ~new_n62_;
  assign new_n64_ = ~new_n63_ | ~new_n17_;
  assign new_n65_ = ~new_n34_;
  assign new_n66_ = ~new_n37_ | ~new_n38_;
  assign new_n67_ = ~x3 & ~x4;
  assign new_n68_ = ~new_n67_ & ~new_n22_;
  assign new_n69_ = ~new_n16_ | ~new_n51_;
  assign new_n70_ = (new_n52_ | new_n69_) & (~new_n33_ | ~new_n29_);
  assign new_n71_ = new_n66_ ? (~new_n68_ ^ new_n70_) : (new_n68_ ^ new_n70_);
  assign new_n72_ = new_n35_ | (~new_n65_ & ~new_n71_);
  assign f4 = ~new_n72_ | ~new_n64_;
  assign f5 = ~new_n46_;
  assign new_n75_ = ~new_n43_ | ~new_n16_;
  assign f6 = new_n75_ & (new_n35_ | new_n54_ | new_n71_);
  assign f7 = ~f8 & (~new_n17_ | ~new_n63_) & (~new_n43_ | ~new_n36_);
  assign f1 = 1'b0;
  assign f9 = new_n75_ & (new_n35_ | new_n54_ | new_n71_);
endmodule


