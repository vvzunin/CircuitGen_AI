module CCGRCG84( x0, x1, x2, x3, f1, f2, f3, f4, f5, f6 );

	input x0, x1, x2, x3;
	output f1, f2, f3, f4, f5, f6;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295;

	nor (d1, x0);
	xnor (d2, x2, x3);
	xnor (d3, x1, x2);
	xnor (d4, x2, x3);
	not (d5, d3);
	and (d6, d1, d2);
	and (d7, d2, d4);
	nor (d8, d2, d4);
	not (d9, d4);
	or (d10, d2, d3);
	and (d11, d4);
	and (d12, d1, d2);
	buf (d13, d4);
	nor (d14, d3, d4);
	nor (d15, d2, d3);
	not (d16, x3);
	or (d17, d2, d4);
	xor (d18, d4);
	xnor (d19, d1, d4);
	not (d20, d1);
	xor (d21, d2, d3);
	buf (d22, d2);
	or (d23, d1, d2);
	xnor (d24, d1, d2);
	and (d25, d2, d3);
	nand (d26, d3, d4);
	not (d27, x0);
	xor (d28, d1, d2);
	or (d29, d1, d3);
	and (d30, d3, d4);
	nand (d31, d3, d4);
	xor (d32, d1, d2);
	or (d33, d2, d4);
	nor (d34, d2, d4);
	or (d35, d2);
	xor (d36, d3);
	nand (d37, d1, d2);
	and (d38, d3, d4);
	buf (d39, x3);
	nand (d40, d1, d3);
	xnor (d41, d3);
	xor (d42, d1);
	and (d43, d3);
	xnor (d44, d2, d3);
	nand (d45, d2, d3);
	nor (d46, d1, d3);
	or (d47, d1, d4);
	nand (d48, d4);
	xnor (d49, d4);
	buf (d50, x2);
	xor (d51, d1, d4);
	and (d52, d1, d3);
	nand (d53, d1);
	nand (d54, d2, d4);
	nor (d55, d3);
	buf (d56, d1);
	xor (d57, d1, d3);
	nand (d58, d1, d3);
	buf (d59, x1);
	and (d60, d2);
	and (d61, d1, d3);
	nor (d62, d1, d2);
	or (d63, d3, d4);
	not (d64, x1);
	and (d65, d2, d4);
	or (d66, d3);
	xor (d67, d2, d4);
	xnor (d68, d7, d21);
	buf (d69, d46);
	nor (d70, d28, d61);
	buf (d71, d26);
	xnor (d72, d24, d50);
	xor (d73, d12, d42);
	and (d74, d20, d52);
	nand (d75, d45, d61);
	not (d76, d64);
	xor (d77, d23, d37);
	nand (d78, d36, d48);
	nand (d79, d43, d59);
	xnor (d80, d12, d65);
	nand (d81, d40, d62);
	and (d82, d7, d61);
	xnor (d83, d34, d60);
	and (d84, d14, d29);
	xor (d85, d58, d61);
	not (d86, d5);
	xnor (d87, d76, d83);
	and (d88, d75, d81);
	xnor (d89, d73, d75);
	or (d90, d80);
	or (d91, d71, d75);
	nand (d92, d73, d82);
	nor (d93, d71, d81);
	xnor (d94, d73, d86);
	nand (d95, d78, d84);
	buf (d96, d68);
	nand (d97, d70, d76);
	xnor (d98, d72, d77);
	buf (d99, d23);
	nor (d100, d75, d85);
	xor (d101, d73, d86);
	nor (d102, d69, d75);
	nand (d103, d68);
	buf (d104, d37);
	nand (d105, d71, d78);
	nor (d106, d70, d74);
	buf (d107, d11);
	nor (d108, d73, d77);
	or (d109, d69, d82);
	and (d110, d69, d75);
	xor (d111, d68, d86);
	xor (d112, d69, d82);
	nor (d113, d76, d80);
	and (d114, d76, d77);
	buf (d115, d75);
	or (d116, d72, d77);
	nand (d117, d70, d76);
	nand (d118, d74, d76);
	xor (d119, d71, d73);
	nor (d120, d71, d84);
	xnor (d121, d71, d82);
	not (d122, d74);
	nor (d123, d78, d84);
	xor (d124, d81, d83);
	xnor (d125, d76, d81);
	xnor (d126, d73, d77);
	xnor (d127, d81, d83);
	xnor (d128, d82, d85);
	xor (d129, d75, d77);
	not (d130, d60);
	and (d131, d70, d77);
	or (d132, d72, d81);
	nor (d133, d77, d83);
	xor (d134, d68, d72);
	nor (d135, d77, d78);
	not (d136, d21);
	xor (d137, d68, d71);
	buf (d138, d51);
	buf (d139, d27);
	xnor (d140, d80, d82);
	and (d141, d68, d80);
	nand (d142, d78, d85);
	or (d143, d82, d86);
	nor (d144, d79, d82);
	and (d145, d73, d84);
	nor (d146, d80, d83);
	or (d147, d68, d80);
	or (d148, d69, d81);
	buf (d149, d20);
	buf (d150, d14);
	xor (d151, d73, d77);
	nand (d152, d75, d86);
	not (d153, d65);
	or (d154, d72, d76);
	and (d155, d75, d77);
	nor (d156, d73, d85);
	and (d157, d79, d80);
	buf (d158, d7);
	xnor (d159, d81, d84);
	nand (d160, d70, d79);
	and (d161, d79, d82);
	nor (d162, d138, d160);
	nand (d163, d106, d113);
	not (d164, d80);
	or (d165, d164);
	nand (d166, d162, d164);
	nor (d167, d162, d164);
	nand (d168, d163);
	xor (d169, d163, d164);
	nor (d170, d163);
	not (d171, d34);
	and (d172, d162, d164);
	buf (d173, d88);
	not (d174, d59);
	xnor (d175, d162, d163);
	and (d176, d162);
	not (d177, d89);
	xor (d178, d162);
	and (d179, d162, d163);
	xor (d180, d163, d164);
	buf (d181, d110);
	buf (d182, d152);
	buf (d183, d57);
	or (d184, d163, d164);
	buf (d185, d81);
	or (d186, d163, d164);
	not (d187, d141);
	nand (d188, d176, d178);
	xnor (d189, d173, d185);
	xor (d190, d171, d187);
	buf (d191, d91);
	xnor (d192, d176, d184);
	nor (d193, d175, d185);
	xnor (d194, d173, d183);
	xor (d195, d177, d186);
	buf (d196, d186);
	xnor (d197, d177, d178);
	or (d198, d179, d180);
	nor (d199, d176, d177);
	nand (d200, d165, d175);
	nand (d201, d171, d186);
	buf (d202, d39);
	not (d203, d163);
	nand (d204, d165, d167);
	not (d205, d35);
	nand (d206, d165, d179);
	or (d207, d170, d177);
	or (d208, d167, d173);
	nor (d209, d176, d181);
	nor (d210, d174, d184);
	not (d211, d36);
	xnor (d212, d166, d169);
	xnor (d213, d167, d176);
	or (d214, d171, d183);
	not (d215, d26);
	xor (d216, d173);
	buf (d217, d17);
	xor (d218, d170, d182);
	xnor (d219, d177);
	xnor (d220, d165, d184);
	nand (d221, d168, d169);
	not (d222, d44);
	not (d223, d133);
	xor (d224, d165, d174);
	nand (d225, d165, d183);
	or (d226, d172, d182);
	xor (d227, d179, d185);
	nor (d228, d175, d180);
	xor (d229, d170, d172);
	xor (d230, d166, d171);
	nor (d231, d178, d180);
	and (d232, d174, d182);
	not (d233, d132);
	and (d234, d182, d187);
	or (d235, d176, d177);
	not (d236, d184);
	buf (d237, d94);
	nor (d238, d181, d185);
	and (d239, d165, d173);
	nand (d240, d176, d185);
	or (d241, d171, d174);
	xor (d242, d172, d184);
	nand (d243, d171, d173);
	not (d244, d29);
	nor (d245, d165, d170);
	and (d246, d167, d177);
	xor (d247, d177, d182);
	and (d248, d165, d169);
	nor (d249, d182);
	nand (d250, d166, d171);
	xor (d251, d174, d183);
	or (d252, d170, d181);
	and (d253, d177, d178);
	or (d254, d182, d187);
	or (d255, d168, d172);
	and (d256, d168, d176);
	and (d257, d178, d184);
	xor (d258, d168, d176);
	nand (d259, d181, d186);
	and (d260, d170, d172);
	or (d261, d165, d182);
	xor (d262, d174, d184);
	nand (d263, d179, d180);
	not (d264, d153);
	nor (d265, d167, d177);
	buf (d266, d84);
	xor (d267, d165, d182);
	nor (d268, d173, d175);
	not (d269, d156);
	xor (d270, d182, d186);
	or (d271, d167, d182);
	nand (d272, d174, d187);
	and (d273, d179, d182);
	nand (d274, d228, d255);
	or (d275, d208, d216);
	nand (d276, d219, d227);
	and (d277, d197, d200);
	xor (d278, d233, d252);
	xnor (d279, d194, d257);
	xnor (d280, d213, d242);
	nor (d281, d223, d273);
	nor (d282, d193, d204);
	or (d283, d216, d254);
	xnor (d284, d257, d271);
	buf (d285, d204);
	buf (d286, d230);
	nor (d287, d197, d218);
	or (d288, d189, d244);
	xnor (d289, d235, d253);
	or (d290, d225, d238);
	or (d291, d190, d225);
	xor (d292, d200, d272);
	xor (d293, d197, d231);
	buf (d294, d143);
	or (d295, d204, d230);
	assign f1 = d277;
	assign f2 = d286;
	assign f3 = d294;
	assign f4 = d288;
	assign f5 = d290;
	assign f6 = d288;
endmodule
