module CCGRCG60( x0, x1, x2, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13 );

	input x0, x1, x2;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159;

	nand (d1, x2);
	nand (d2, x1, x2);
	not (d3, x0);
	buf (d4, x2);
	and (d5, x0, x2);
	xnor (d6, x2);
	nand (d7, x0);
	xnor (d8, x0, x2);
	not (d9, x1);
	buf (d10, x1);
	and (d11, x2);
	xnor (d12, x0, x2);
	not (d13, x2);
	xor (d14, x2);
	nor (d15, x0, x1);
	xor (d16, x1, x2);
	or (d17, x2);
	or (d18, x0, x1);
	nor (d19, x2);
	nor (d20, x0, x2);
	and (d21, x0);
	and (d22, x0, x1);
	and (d23, x1, x2);
	nor (d24, x0, x2);
	xnor (d25, x1, x2);
	nand (d26, x1, x2);
	or (d27, x1);
	and (d28, x0, x1);
	xor (d29, x0, x1);
	xor (d30, x0, x2);
	nor (d31, x1, x2);
	buf (d32, x0);
	or (d33, x1, x2);
	or (d34, x0, x1);
	xnor (d35, x0, x1);
	xor (d36, x0);
	nor (d37, x1, x2);
	and (d38, x1);
	nand (d39, x0, x1);
	or (d40, x0, x2);
	nor (d41, x1);
	nand (d42, x0, x2);
	nor (d43, x0, x1);
	xnor (d44, x1);
	nor (d45, x0);
	or (d46, d13, d41);
	xnor (d47, d17, d36);
	nand (d48, d8, d18);
	buf (d49, d32);
	buf (d50, d22);
	and (d51, d42, d44);
	nand (d52, d14, d22);
	xor (d53, d5, d16);
	or (d54, d5, d9);
	or (d55, d6, d28);
	nand (d56, d8, d31);
	xor (d57, d16, d24);
	or (d58, d13, d32);
	and (d59, d14, d40);
	nand (d60, d5, d45);
	buf (d61, d1);
	nand (d62, d7, d22);
	and (d63, d23, d31);
	nand (d64, d19, d43);
	buf (d65, d18);
	nor (d66, d5, d42);
	or (d67, d1, d29);
	and (d68, d46, d62);
	buf (d69, d25);
	not (d70, d16);
	nand (d71, d51, d67);
	xnor (d72, d49, d60);
	and (d73, d54, d62);
	nand (d74, d55, d66);
	not (d75, d19);
	and (d76, d49, d65);
	not (d77, d2);
	xor (d78, d48, d63);
	nor (d79, d57, d60);
	and (d80, d57, d61);
	xnor (d81, d54, d67);
	nor (d82, d49);
	nor (d83, d59, d65);
	buf (d84, d36);
	xor (d85, d60, d65);
	xnor (d86, d50, d56);
	not (d87, d51);
	buf (d88, d11);
	nand (d89, d56, d57);
	not (d90, d66);
	not (d91, d57);
	nand (d92, d53, d54);
	nand (d93, d49, d54);
	xnor (d94, d48, d59);
	or (d95, d64, d67);
	xor (d96, d60, d64);
	xor (d97, d57, d65);
	not (d98, d40);
	nor (d99, d55, d60);
	xor (d100, d47, d64);
	nand (d101, d57, d67);
	not (d102, d9);
	nand (d103, d52, d60);
	nor (d104, d46, d53);
	and (d105, d46, d50);
	not (d106, d29);
	nand (d107, d57, d64);
	and (d108, d57, d66);
	nand (d109, d58, d61);
	nor (d110, d56, d66);
	buf (d111, d51);
	xor (d112, d64);
	nor (d113, d48, d52);
	nor (d114, d46, d59);
	nand (d115, d62, d67);
	nand (d116, d49, d58);
	and (d117, d46, d66);
	and (d118, d54, d57);
	or (d119, d56, d58);
	or (d120, d48, d64);
	not (d121, d33);
	nand (d122, d63, d64);
	xnor (d123, d55, d57);
	or (d124, d55, d62);
	and (d125, d46, d50);
	buf (d126, d12);
	nand (d127, d59, d67);
	not (d128, d20);
	xor (d129, d48, d52);
	xnor (d130, d50, d55);
	buf (d131, d31);
	and (d132, d57, d62);
	xor (d133, d58, d59);
	or (d134, d51, d56);
	not (d135, d67);
	nor (d136, d51, d67);
	or (d137, d54, d65);
	xor (d138, d48, d65);
	and (d139, d60);
	buf (d140, d137);
	and (d141, d90, d102);
	xor (d142, d108, d115);
	xnor (d143, d117, d138);
	xnor (d144, d132, d139);
	not (d145, d86);
	nor (d146, d100, d128);
	xor (d147, d101, d126);
	not (d148, d5);
	not (d149, d73);
	nor (d150, d80, d110);
	not (d151, d90);
	xor (d152, d81, d91);
	or (d153, d72, d110);
	and (d154, d104, d113);
	nand (d155, d93, d124);
	not (d156, d101);
	nor (d157, d75, d131);
	buf (d158, d71);
	buf (d159, d14);
	assign f1 = d149;
	assign f2 = d148;
	assign f3 = d159;
	assign f4 = d153;
	assign f5 = d157;
	assign f6 = d150;
	assign f7 = d147;
	assign f8 = d152;
	assign f9 = d141;
	assign f10 = d149;
	assign f11 = d143;
	assign f12 = d156;
	assign f13 = d148;
endmodule
