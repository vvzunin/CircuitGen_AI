module CCGRCG166( x0, x1, x2, x3, x4, x5, f1, f2, f3, f4, f5, f6, f7, f8, f9 );

	input x0, x1, x2, x3, x4, x5;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314, d315, d316, d317, d318, d319, d320, d321, d322, d323, d324, d325, d326, d327, d328, d329, d330, d331, d332, d333, d334, d335, d336, d337, d338, d339, d340, d341, d342, d343, d344, d345, d346, d347, d348, d349, d350, d351, d352, d353, d354, d355, d356, d357, d358, d359, d360, d361, d362, d363, d364, d365;

	nor (d1, x4, x5);
	nand (d2, x3, x4);
	buf (d3, x4);
	buf (d4, x0);
	and (d5, x0, x3);
	or (d6, x1, x3);
	xnor (d7, x0, x1);
	xnor (d8, x4, x5);
	and (d9, x0, x2);
	or (d10, d6, d7);
	buf (d11, d2);
	buf (d12, d8);
	or (d13, d1, d5);
	xnor (d14, d6, d8);
	nand (d15, d1, d9);
	and (d16, d4, d6);
	xnor (d17, d3, d5);
	nor (d18, d1, d5);
	nand (d19, d10, d13);
	or (d20, d14, d17);
	not (d21, d7);
	xnor (d22, d12, d16);
	not (d23, x1);
	and (d24, d12, d18);
	or (d25, d12, d13);
	xor (d26, d11, d15);
	nor (d27, d13, d15);
	xor (d28, d10, d13);
	xnor (d29, d15, d17);
	or (d30, d12, d13);
	xor (d31, d10, d18);
	xnor (d32, d14, d15);
	buf (d33, d13);
	not (d34, d5);
	xnor (d35, d12, d15);
	xnor (d36, d11, d18);
	or (d37, d13, d15);
	or (d38, d11);
	nand (d39, d14, d18);
	xor (d40, d12, d18);
	and (d41, d10, d14);
	nand (d42, d14, d18);
	not (d43, d17);
	nand (d44, d12, d15);
	xnor (d45, d10, d13);
	xor (d46, d11, d14);
	or (d47, d12, d16);
	xor (d48, d12, d14);
	nor (d49, d11, d17);
	not (d50, d9);
	buf (d51, d18);
	not (d52, d1);
	not (d53, x4);
	and (d54, d15);
	nor (d55, d11, d12);
	xor (d56, d13, d14);
	and (d57, d15, d16);
	xor (d58, d17, d18);
	not (d59, x2);
	buf (d60, d10);
	xor (d61, d15);
	or (d62, d10, d16);
	or (d63, d16);
	xor (d64, d15, d17);
	or (d65, d15, d18);
	nor (d66, d13, d14);
	nand (d67, d13, d16);
	or (d68, d16, d18);
	or (d69, d13, d17);
	buf (d70, d17);
	xor (d71, d12, d15);
	and (d72, d10, d15);
	xnor (d73, d11, d12);
	xor (d74, d14);
	nor (d75, d12, d14);
	not (d76, d36);
	xor (d77, d65, d72);
	xnor (d78, d41, d61);
	and (d79, d42, d72);
	or (d80, d58, d66);
	not (d81, d21);
	buf (d82, d72);
	not (d83, x5);
	xnor (d84, d54, d64);
	buf (d85, d31);
	nand (d86, d24, d40);
	or (d87, d37, d49);
	or (d88, d36, d50);
	xor (d89, d29, d38);
	xnor (d90, d28, d59);
	xnor (d91, d28, d72);
	buf (d92, d69);
	and (d93, d43, d68);
	nor (d94, d49, d74);
	xor (d95, d37, d66);
	and (d96, d26, d37);
	or (d97, d27, d35);
	nand (d98, d51, d58);
	xor (d99, d21, d32);
	xor (d100, d22, d44);
	buf (d101, d16);
	and (d102, d34, d60);
	not (d103, d11);
	nor (d104, d59, d73);
	xor (d105, d29, d56);
	xor (d106, d31, d54);
	or (d107, d36, d67);
	xnor (d108, d42, d44);
	xor (d109, d44, d66);
	and (d110, d37, d39);
	or (d111, d37, d53);
	xor (d112, d21, d35);
	nand (d113, d52, d72);
	or (d114, d45, d59);
	nand (d115, d28, d29);
	not (d116, d74);
	buf (d117, d52);
	nand (d118, d43, d74);
	buf (d119, d19);
	nor (d120, d20, d37);
	and (d121, d95, d110);
	not (d122, d99);
	or (d123, d89, d117);
	xor (d124, d78, d95);
	nor (d125, d83, d90);
	and (d126, d85, d102);
	xnor (d127, d78, d117);
	xor (d128, d96, d97);
	xor (d129, d81, d88);
	not (d130, d52);
	or (d131, d104, d108);
	and (d132, d87, d94);
	xnor (d133, d82, d116);
	and (d134, d109, d113);
	not (d135, d46);
	or (d136, d102, d103);
	and (d137, d76, d89);
	buf (d138, d90);
	or (d139, d102, d115);
	and (d140, d80, d84);
	xnor (d141, d85, d93);
	xor (d142, d82, d113);
	buf (d143, d5);
	buf (d144, d40);
	buf (d145, d55);
	xor (d146, d84, d99);
	xnor (d147, d90, d118);
	or (d148, d79, d88);
	xor (d149, d84, d92);
	nand (d150, d109, d110);
	and (d151, d111, d118);
	or (d152, d77, d111);
	xor (d153, d94, d110);
	nor (d154, d78, d103);
	nand (d155, d81, d100);
	xnor (d156, d93, d96);
	xnor (d157, d108, d116);
	not (d158, d35);
	buf (d159, d92);
	or (d160, d90, d110);
	nand (d161, d78, d109);
	xor (d162, d77, d115);
	not (d163, d30);
	xor (d164, d94, d104);
	buf (d165, d33);
	nand (d166, d93, d111);
	or (d167, d93, d107);
	and (d168, d83, d91);
	not (d169, d80);
	xor (d170, d76, d96);
	xor (d171, d94, d109);
	xnor (d172, d109, d115);
	not (d173, d58);
	xor (d174, d90, d104);
	or (d175, d123, d155);
	xor (d176, d153, d154);
	buf (d177, d143);
	xnor (d178, d139, d159);
	nor (d179, d133, d163);
	xor (d180, d134, d136);
	and (d181, d122, d159);
	buf (d182, d141);
	not (d183, d23);
	xor (d184, d144);
	not (d185, d101);
	or (d186, d124, d143);
	nand (d187, d124, d174);
	xnor (d188, d130, d169);
	xor (d189, d136, d157);
	not (d190, d124);
	or (d191, d146, d157);
	nor (d192, d127, d172);
	xnor (d193, d135, d170);
	or (d194, d135, d157);
	nand (d195, d125, d145);
	nand (d196, d126, d132);
	and (d197, d142, d173);
	not (d198, d29);
	xor (d199, d160, d166);
	or (d200, d147, d157);
	or (d201, d186, d200);
	or (d202, d186, d188);
	buf (d203, d62);
	and (d204, d181, d196);
	xnor (d205, d182, d185);
	xor (d206, d187, d197);
	and (d207, d182, d187);
	and (d208, d186, d187);
	and (d209, d189, d194);
	and (d210, d196, d197);
	xor (d211, d179, d200);
	or (d212, d179, d200);
	not (d213, d60);
	xor (d214, d175, d188);
	and (d215, d182, d183);
	and (d216, d176, d191);
	and (d217, d190, d191);
	xnor (d218, d181, d191);
	or (d219, d177, d182);
	nor (d220, d186, d189);
	nand (d221, d177, d198);
	not (d222, d194);
	buf (d223, d125);
	xnor (d224, d181, d197);
	nor (d225, d182, d194);
	buf (d226, d163);
	and (d227, d197);
	nor (d228, d179, d188);
	nor (d229, d185, d197);
	buf (d230, d7);
	xnor (d231, d179, d183);
	or (d232, d178, d183);
	buf (d233, d193);
	buf (d234, d175);
	not (d235, d34);
	buf (d236, d166);
	nand (d237, d175, d188);
	nand (d238, d185, d199);
	and (d239, d180, d185);
	nor (d240, d195);
	xor (d241, d176, d183);
	buf (d242, d172);
	buf (d243, d196);
	xnor (d244, d192, d196);
	nor (d245, d186, d198);
	buf (d246, d183);
	nor (d247, d182, d185);
	not (d248, d4);
	or (d249, d182, d197);
	buf (d250, d162);
	xnor (d251, d177, d192);
	and (d252, d179, d198);
	or (d253, d187, d197);
	nand (d254, d185, d193);
	nand (d255, d176, d198);
	xor (d256, d192, d193);
	nand (d257, d176, d178);
	not (d258, d69);
	xnor (d259, d186, d197);
	nand (d260, d180, d186);
	not (d261, d70);
	not (d262, d120);
	nor (d263, d184, d193);
	nand (d264, d179, d199);
	xor (d265, d188, d196);
	buf (d266, d32);
	nor (d267, d175, d192);
	not (d268, d44);
	nor (d269, d176, d186);
	nand (d270, d182, d190);
	nand (d271, d182, d188);
	buf (d272, d86);
	xnor (d273, d186, d188);
	not (d274, d43);
	not (d275, d131);
	buf (d276, d63);
	xor (d277, d183, d193);
	nor (d278, d184, d195);
	xor (d279, d185, d188);
	xnor (d280, d186, d192);
	nor (d281, d180, d195);
	xor (d282, d192, d198);
	buf (d283, d82);
	not (d284, d67);
	nand (d285, d191, d195);
	and (d286, d185, d196);
	xor (d287, d186, d191);
	buf (d288, d87);
	and (d289, d179, d185);
	xnor (d290, d193, d198);
	nand (d291, d176, d189);
	or (d292, d237, d274);
	xor (d293, d247, d263);
	nand (d294, d215, d234);
	buf (d295, d153);
	not (d296, d168);
	nand (d297, d221, d236);
	xnor (d298, d214, d248);
	nand (d299, d232, d247);
	nand (d300, d220, d271);
	or (d301, d207, d259);
	xor (d302, d218, d239);
	not (d303, d155);
	nand (d304, d206, d227);
	xnor (d305, d246, d289);
	xnor (d306, d233, d247);
	nand (d307, d216, d217);
	xnor (d308, d220, d226);
	xnor (d309, d246, d282);
	buf (d310, d230);
	or (d311, d201, d204);
	and (d312, d211, d254);
	nor (d313, d231, d253);
	and (d314, d232, d282);
	or (d315, d265, d284);
	and (d316, d217, d222);
	or (d317, d222, d284);
	xor (d318, d201, d279);
	nand (d319, d225, d278);
	not (d320, d144);
	not (d321, d251);
	nand (d322, d300, d311);
	not (d323, d91);
	not (d324, d264);
	buf (d325, d160);
	buf (d326, d219);
	and (d327, d302, d313);
	buf (d328, d57);
	or (d329, d314, d316);
	xor (d330, d297, d301);
	or (d331, d302, d308);
	buf (d332, d103);
	buf (d333, d173);
	xnor (d334, d294, d298);
	or (d335, d296, d297);
	nand (d336, d301, d317);
	and (d337, d309, d315);
	and (d338, d299, d317);
	or (d339, d293, d316);
	buf (d340, d30);
	not (d341, d262);
	or (d342, d308, d319);
	nor (d343, d293, d297);
	and (d344, d301);
	buf (d345, d12);
	xnor (d346, d338, d341);
	buf (d347, d269);
	or (d348, d327, d343);
	nand (d349, d335);
	nand (d350, d339, d344);
	and (d351, d327, d328);
	and (d352, d323, d336);
	or (d353, d321, d333);
	nand (d354, d324, d345);
	and (d355, d330, d336);
	nand (d356, d323, d345);
	nand (d357, d326, d342);
	and (d358, d327, d331);
	nor (d359, d328, d332);
	or (d360, d326, d331);
	not (d361, d309);
	xnor (d362, d326, d336);
	and (d363, d333, d345);
	xor (d364, d323, d326);
	buf (d365, d277);
	assign f1 = d361;
	assign f2 = d362;
	assign f3 = d362;
	assign f4 = d347;
	assign f5 = d363;
	assign f6 = d346;
	assign f7 = d365;
	assign f8 = d348;
	assign f9 = d358;
endmodule
