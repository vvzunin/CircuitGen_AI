module CCGRCG165( x0, x1, x2, x3, x4, x5, f1, f2, f3, f4, f5, f6, f7, f8 );

	input x0, x1, x2, x3, x4, x5;
	output f1, f2, f3, f4, f5, f6, f7, f8;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41;

	or (d1, x0, x5);
	or (d2, x1, x5);
	xor (d3, x0, x1);
	buf (d4, x0);
	nor (d5, x0, x3);
	nor (d6, x0, x1);
	or (d7, x0, x4);
	and (d8, x4);
	xnor (d9, x2, x5);
	buf (d10, x2);
	xnor (d11, x0, x3);
	xor (d12, x0, x4);
	or (d13, x1, x3);
	nand (d14, x0, x4);
	nor (d15, x3, x4);
	nor (d16, x1, x5);
	xor (d17, x5);
	nor (d18, x0, x4);
	buf (d19, x5);
	buf (d20, x4);
	not (d21, x2);
	not (d22, x3);
	nand (d23, x3);
	xor (d24, x3, x5);
	and (d25, x0, x5);
	or (d26, x1, x4);
	nor (d27, x2, x4);
	nor (d28, x2, x5);
	or (d29, x1, x2);
	and (d30, x0, x4);
	nor (d31, x1, x3);
	nor (d32, x4, x5);
	buf (d33, x1);
	xor (d34, x0, x2);
	xnor (d35, x1, x3);
	xnor (d36, x4, x5);
	or (d37, x0, x3);
	xor (d38, x0);
	and (d39, x2, x5);
	nand (d40, x0, x1);
	and (d41, x0, x2);
	assign f1 = d3;
	assign f2 = d14;
	assign f3 = d12;
	assign f4 = d25;
	assign f5 = d19;
	assign f6 = d24;
	assign f7 = d4;
	assign f8 = d28;
endmodule
