module CCGRCG151( x0, x1, x2, x3, x4, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17, f18, f19, f20 );

	input x0, x1, x2, x3, x4;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17, f18, f19, f20;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314, d315, d316, d317, d318, d319, d320, d321, d322, d323, d324, d325, d326, d327, d328, d329, d330, d331, d332, d333, d334, d335, d336, d337, d338, d339, d340, d341, d342, d343, d344, d345, d346, d347, d348, d349, d350, d351, d352, d353, d354, d355, d356, d357, d358, d359, d360, d361, d362, d363, d364, d365, d366, d367, d368, d369, d370, d371, d372, d373, d374, d375, d376, d377, d378, d379, d380, d381, d382, d383, d384, d385, d386, d387, d388, d389, d390, d391, d392, d393, d394, d395, d396, d397, d398, d399, d400, d401, d402, d403, d404, d405, d406, d407, d408, d409, d410, d411, d412, d413, d414, d415, d416, d417, d418, d419, d420, d421, d422, d423, d424, d425, d426, d427, d428, d429, d430, d431, d432, d433, d434, d435;

	nor (d1, x1, x2);
	buf (d2, x0);
	nand (d3, x1, x3);
	nor (d4, x3, x4);
	nand (d5, x2, x4);
	not (d6, x0);
	xor (d7, x1, x3);
	and (d8, x3, x4);
	nor (d9, x1, x4);
	buf (d10, x4);
	or (d11, x1, x2);
	nand (d12, x0, x4);
	nand (d13, x0, x2);
	xor (d14, x1, x4);
	or (d15, x0, x3);
	buf (d16, x3);
	nor (d17, x0, x1);
	and (d18, x1, x2);
	nand (d19, x2, x4);
	or (d20, x0, x4);
	xor (d21, x2);
	and (d22, x1, x2);
	xnor (d23, x0, x1);
	not (d24, x2);
	nor (d25, x0, x2);
	or (d26, x0, x3);
	nor (d27, x2, x4);
	and (d28, x3);
	nand (d29, x3, x4);
	nor (d30, x1, x3);
	nor (d31, x0);
	or (d32, x4);
	nand (d33, x0, x1);
	not (d34, x4);
	xor (d35, x1, x4);
	or (d36, x1, x4);
	or (d37, x3, x4);
	or (d38, x2, x4);
	or (d39, x2, x3);
	xnor (d40, x3, x4);
	xnor (d41, x0, x3);
	or (d42, x0);
	nor (d43, x2, x4);
	nand (d44, x1, x2);
	and (d45, x2, x3);
	and (d46, x3, x4);
	xnor (d47, x0, x3);
	xor (d48, x1, x2);
	buf (d49, x2);
	or (d50, x0, x1);
	xor (d51, x1, x2);
	nor (d52, x0, x2);
	nor (d53, x1, x3);
	nor (d54, x0, x3);
	nor (d55, x0, x4);
	not (d56, d44);
	or (d57, d5, d24);
	buf (d58, d16);
	not (d59, d39);
	not (d60, d36);
	and (d61, d37, d42);
	not (d62, d14);
	nand (d63, d32, d41);
	buf (d64, x1);
	nand (d65, d27, d54);
	xnor (d66, d3, d50);
	nor (d67, d46, d47);
	xor (d68, d1, d14);
	xor (d69, d22, d55);
	nand (d70, d17, d41);
	nand (d71, d4, d14);
	not (d72, d32);
	nand (d73, d19, d34);
	xnor (d74, d11, d23);
	not (d75, d22);
	not (d76, d31);
	nand (d77, d36, d55);
	nand (d78, d42, d55);
	buf (d79, d41);
	nor (d80, d35, d45);
	nand (d81, d19, d44);
	nor (d82, d10, d49);
	and (d83, d26, d31);
	nand (d84, d27, d39);
	or (d85, d57, d67);
	xor (d86, d63, d77);
	xor (d87, d77, d81);
	and (d88, d59, d69);
	xor (d89, d75, d81);
	not (d90, d42);
	or (d91, d76, d79);
	xor (d92, d70, d81);
	nor (d93, d72, d75);
	xor (d94, d67, d84);
	xnor (d95, d57, d72);
	nand (d96, d81, d82);
	buf (d97, d34);
	not (d98, d34);
	xnor (d99, d63, d84);
	and (d100, d63, d64);
	nand (d101, d69, d79);
	nand (d102, d75, d77);
	and (d103, d56, d67);
	nor (d104, d66, d80);
	buf (d105, d75);
	or (d106, d64, d80);
	not (d107, d78);
	xor (d108, d62, d67);
	xor (d109, d69, d79);
	nand (d110, d58, d73);
	xnor (d111, d78, d79);
	nor (d112, d62, d83);
	nand (d113, d77, d78);
	or (d114, d68, d70);
	nor (d115, d60, d61);
	nor (d116, d60, d76);
	buf (d117, d6);
	nor (d118, d61, d80);
	nand (d119, d67, d78);
	or (d120, d71, d73);
	nor (d121, d63, d76);
	nor (d122, d68, d83);
	nand (d123, d74, d80);
	xor (d124, d79, d81);
	buf (d125, d79);
	xor (d126, d62, d74);
	nor (d127, d59, d79);
	xnor (d128, d68, d70);
	or (d129, d66, d77);
	nor (d130, d79, d80);
	buf (d131, d1);
	buf (d132, d47);
	xor (d133, d62, d83);
	and (d134, d76, d83);
	and (d135, d73, d75);
	not (d136, d82);
	not (d137, d64);
	buf (d138, d60);
	or (d139, d134, d135);
	not (d140, d67);
	xnor (d141, d111, d128);
	xor (d142, d118, d129);
	or (d143, d90, d111);
	nand (d144, d93, d112);
	xnor (d145, d101, d108);
	or (d146, d97, d101);
	nand (d147, d118, d120);
	xor (d148, d126, d135);
	xor (d149, d90, d104);
	nor (d150, d117, d130);
	or (d151, d120, d126);
	nand (d152, d89, d90);
	nor (d153, d89, d101);
	xor (d154, d112, d126);
	xnor (d155, d91, d101);
	not (d156, d70);
	buf (d157, d61);
	nand (d158, d90, d98);
	or (d159, d89, d103);
	nand (d160, d91, d111);
	nor (d161, d86, d100);
	xnor (d162, d121, d129);
	or (d163, d89, d127);
	xor (d164, d94, d125);
	xor (d165, d117, d128);
	and (d166, d94, d108);
	and (d167, d85, d100);
	not (d168, d89);
	xnor (d169, d109);
	buf (d170, d110);
	xnor (d171, d102, d105);
	and (d172, d121, d135);
	and (d173, d96, d98);
	nor (d174, d98, d129);
	nand (d175, d114, d127);
	and (d176, d103, d124);
	and (d177, d93, d126);
	not (d178, d84);
	xor (d179, d102, d116);
	not (d180, d72);
	xnor (d181, d124, d128);
	not (d182, d47);
	nand (d183, d89, d121);
	xnor (d184, d96, d121);
	nand (d185, d87, d124);
	nand (d186, d99, d102);
	not (d187, d21);
	and (d188, d87, d118);
	xor (d189, d93, d130);
	not (d190, d76);
	not (d191, d129);
	nor (d192, d95, d100);
	not (d193, d122);
	nor (d194, d124, d128);
	buf (d195, d63);
	and (d196, d96, d122);
	xnor (d197, d108, d115);
	not (d198, d93);
	buf (d199, d43);
	nand (d200, d99, d133);
	xnor (d201, d120, d124);
	xor (d202, d119, d120);
	or (d203, d98, d118);
	and (d204, d96, d107);
	xnor (d205, d100, d133);
	not (d206, d88);
	nor (d207, d89, d100);
	not (d208, d16);
	or (d209, d96, d131);
	buf (d210, d122);
	xor (d211, d86, d116);
	and (d212, d101, d132);
	not (d213, d130);
	buf (d214, d128);
	not (d215, d112);
	and (d216, d121, d132);
	not (d217, d79);
	or (d218, d110, d127);
	or (d219, d86, d107);
	buf (d220, d80);
	nand (d221, d108, d120);
	and (d222, d108, d126);
	xnor (d223, d94, d121);
	buf (d224, d56);
	xnor (d225, d107, d109);
	and (d226, d110, d121);
	not (d227, d54);
	not (d228, d4);
	or (d229, d129, d131);
	xor (d230, d94, d113);
	and (d231, d90, d124);
	buf (d232, d57);
	not (d233, d116);
	buf (d234, d88);
	nand (d235, d197, d200);
	buf (d236, d226);
	buf (d237, d217);
	nand (d238, d190, d214);
	not (d239, d138);
	nand (d240, d138, d207);
	nor (d241, d141, d169);
	xor (d242, d197, d210);
	not (d243, d20);
	nand (d244, d143, d211);
	nor (d245, d143, d201);
	nand (d246, d145, d192);
	xor (d247, d202, d207);
	buf (d248, d72);
	or (d249, d182, d230);
	nor (d250, d150, d198);
	buf (d251, d197);
	buf (d252, d111);
	xor (d253, d196, d208);
	and (d254, d187, d220);
	xnor (d255, d207, d214);
	and (d256, d148, d222);
	buf (d257, d150);
	xnor (d258, d167, d225);
	not (d259, d226);
	not (d260, d101);
	nor (d261, d137, d156);
	buf (d262, d121);
	xor (d263, d168, d217);
	or (d264, d180, d200);
	xnor (d265, d151, d177);
	or (d266, d182, d222);
	and (d267, d155, d224);
	not (d268, d115);
	or (d269, d153, d165);
	or (d270, d138, d164);
	or (d271, d197, d200);
	or (d272, d148, d219);
	xor (d273, d162, d196);
	and (d274, d198, d204);
	not (d275, d29);
	xor (d276, d169, d176);
	buf (d277, d167);
	not (d278, d157);
	not (d279, d96);
	xor (d280, d203, d228);
	nor (d281, d252, d272);
	xor (d282, d262, d269);
	and (d283, d241, d276);
	buf (d284, d24);
	nor (d285, d255, d275);
	and (d286, d234, d248);
	xnor (d287, d239, d245);
	xnor (d288, d235, d262);
	nand (d289, d241, d279);
	nor (d290, d267, d269);
	xor (d291, d247, d279);
	xnor (d292, d276, d280);
	nand (d293, d258, d278);
	not (d294, d18);
	and (d295, d252, d266);
	not (d296, d25);
	xnor (d297, d277, d278);
	nand (d298, d235, d237);
	or (d299, d245, d260);
	xor (d300, d233, d244);
	xor (d301, d273, d278);
	or (d302, d234, d279);
	xnor (d303, d236, d254);
	xnor (d304, d241, d251);
	xnor (d305, d234, d272);
	and (d306, d260, d279);
	or (d307, d238, d261);
	not (d308, d272);
	not (d309, d212);
	nand (d310, d239, d279);
	nand (d311, d244, d249);
	nand (d312, d265, d275);
	xor (d313, d255, d266);
	or (d314, d238, d250);
	xnor (d315, d246, d254);
	nand (d316, d246, d274);
	buf (d317, d228);
	and (d318, d238, d270);
	nor (d319, d246, d258);
	nand (d320, d241, d268);
	xnor (d321, d237, d271);
	buf (d322, d231);
	xor (d323, d262, d267);
	xor (d324, d237, d242);
	not (d325, d234);
	or (d326, d274, d280);
	and (d327, d238, d268);
	buf (d328, d100);
	or (d329, d265, d275);
	or (d330, d241, d248);
	or (d331, d258, d270);
	xnor (d332, d233, d278);
	nor (d333, d234, d279);
	nor (d334, d257, d270);
	or (d335, d234, d242);
	xor (d336, d246, d253);
	xor (d337, d235, d272);
	not (d338, d139);
	and (d339, d237, d249);
	nor (d340, d286, d337);
	nand (d341, d300, d310);
	xor (d342, d286, d294);
	not (d343, d169);
	buf (d344, d85);
	not (d345, d279);
	xor (d346, d289, d294);
	and (d347, d286, d293);
	buf (d348, d146);
	nand (d349, d317, d337);
	nor (d350, d298, d313);
	nor (d351, d299, d338);
	buf (d352, d2);
	nor (d353, d284, d287);
	nor (d354, d309, d327);
	buf (d355, d254);
	or (d356, d313, d325);
	not (d357, d250);
	nor (d358, d285, d288);
	and (d359, d328, d331);
	or (d360, d284, d321);
	xnor (d361, d323, d326);
	buf (d362, d267);
	nand (d363, d312, d316);
	xor (d364, d299, d331);
	or (d365, d312, d333);
	nand (d366, d298, d317);
	xor (d367, d338);
	nor (d368, d319, d330);
	nor (d369, d292, d320);
	nand (d370, d295, d326);
	nand (d371, d305, d334);
	nand (d372, d290, d333);
	nor (d373, d284, d330);
	nor (d374, d293, d306);
	or (d375, d317, d333);
	not (d376, d98);
	xnor (d377, d349, d371);
	or (d378, d357, d363);
	nor (d379, d363, d369);
	buf (d380, d331);
	xnor (d381, d344, d355);
	or (d382, d362, d369);
	or (d383, d357, d373);
	or (d384, d350, d364);
	or (d385, d352, d356);
	xor (d386, d361, d362);
	xor (d387, d341, d361);
	nor (d388, d340, d346);
	and (d389, d343, d370);
	or (d390, d346, d355);
	or (d391, d351, d359);
	xor (d392, d352, d373);
	and (d393, d344, d365);
	or (d394, d355, d365);
	xor (d395, d340, d350);
	or (d396, d344, d365);
	or (d397, d355, d370);
	nor (d398, d343, d349);
	or (d399, d345, d359);
	buf (d400, d50);
	and (d401, d348, d368);
	buf (d402, d351);
	buf (d403, d89);
	and (d404, d341, d368);
	and (d405, d368);
	not (d406, d66);
	and (d407, d341, d360);
	or (d408, d360, d365);
	xnor (d409, d362, d375);
	or (d410, d370, d374);
	xor (d411, d343, d354);
	xnor (d412, d368, d375);
	xnor (d413, d343, d349);
	xnor (d414, d363, d372);
	and (d415, d365, d369);
	xnor (d416, d357, d369);
	xor (d417, d352, d362);
	not (d418, d266);
	and (d419, d358, d360);
	buf (d420, d342);
	xnor (d421, d361, d370);
	and (d422, d345, d372);
	or (d423, d361, d374);
	buf (d424, d302);
	and (d425, d341, d367);
	xnor (d426, d352, d372);
	xor (d427, d359, d364);
	or (d428, d371, d372);
	nor (d429, d342, d345);
	xnor (d430, d342, d359);
	or (d431, d356, d369);
	not (d432, d189);
	buf (d433, d202);
	xor (d434, d344, d361);
	not (d435, d366);
	assign f1 = d430;
	assign f2 = d385;
	assign f3 = d397;
	assign f4 = d427;
	assign f5 = d382;
	assign f6 = d391;
	assign f7 = d384;
	assign f8 = d403;
	assign f9 = d418;
	assign f10 = d386;
	assign f11 = d416;
	assign f12 = d387;
	assign f13 = d377;
	assign f14 = d400;
	assign f15 = d403;
	assign f16 = d429;
	assign f17 = d423;
	assign f18 = d411;
	assign f19 = d389;
	assign f20 = d402;
endmodule
