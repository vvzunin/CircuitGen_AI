module CCGRCG74( x0, x1, x2, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17, f18, f19, f20 );

	input x0, x1, x2;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17, f18, f19, f20;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120;

	nand (d1, x1, x2);
	or (d2, x0, x2);
	xnor (d3, x1, x2);
	nand (d4, x0);
	and (d5, x1, x2);
	nand (d6, x1, x2);
	nor (d7, x0, x1);
	nor (d8, x1, x2);
	buf (d9, x2);
	not (d10, x1);
	xor (d11, x1, x2);
	xnor (d12, x0, x2);
	not (d13, x0);
	or (d14, x1, x2);
	xor (d15, x0, x1);
	nor (d16, x0);
	nand (d17, x2);
	and (d18, x1, x2);
	nand (d19, x0, x1);
	nand (d20, x0, x1);
	or (d21, x0, x1);
	buf (d22, x1);
	buf (d23, x0);
	not (d24, x2);
	or (d25, x0);
	xnor (d26, x2);
	xor (d27, x1);
	nor (d28, x1, x2);
	xor (d29, x0, x2);
	or (d30, x1, x2);
	xnor (d31, x1, x2);
	xor (d32, x2);
	nand (d33, x0, x2);
	or (d34, x0, x2);
	and (d35, x0, x1);
	xor (d36, x1, x2);
	nor (d37, x0, x1);
	and (d38, x0, x2);
	and (d39, x0, x1);
	xnor (d40, x0);
	nand (d41, d2, d7);
	and (d42, d5, d9);
	or (d43, d4, d36);
	not (d44, d26);
	nor (d45, d42);
	nand (d46, d41, d44);
	nor (d47, d41);
	xnor (d48, d42, d44);
	xor (d49, d44);
	nand (d50, d43, d44);
	nor (d51, d42, d44);
	xor (d52, d41, d42);
	not (d53, d36);
	buf (d54, d15);
	or (d55, d42, d44);
	not (d56, d18);
	nor (d57, d44);
	nor (d58, d43, d44);
	xor (d59, d43, d44);
	or (d60, d41, d43);
	nand (d61, d43, d44);
	nand (d62, d43);
	or (d63, d42, d44);
	and (d64, d41, d43);
	and (d65, d41, d44);
	xor (d66, d41);
	not (d67, d4);
	or (d68, d41, d44);
	nor (d69, d41, d43);
	and (d70, d41, d42);
	nand (d71, d42, d44);
	not (d72, d21);
	buf (d73, d2);
	not (d74, d29);
	not (d75, d41);
	buf (d76, d6);
	or (d77, d43, d44);
	buf (d78, d7);
	and (d79, d55, d67);
	and (d80, d48, d70);
	buf (d81, d59);
	not (d82, d64);
	buf (d83, d1);
	not (d84, d66);
	or (d85, d69, d75);
	nor (d86, d52, d62);
	buf (d87, d27);
	buf (d88, d44);
	xor (d89, d49, d60);
	not (d90, d11);
	nor (d91, d62, d71);
	and (d92, d54, d65);
	and (d93, d50, d76);
	nor (d94, d56, d58);
	buf (d95, d73);
	xnor (d96, d62, d72);
	or (d97, d46, d62);
	not (d98, d35);
	xor (d99, d51, d65);
	xor (d100, d49, d50);
	buf (d101, d20);
	and (d102, d45, d57);
	nand (d103, d46, d54);
	or (d104, d66, d67);
	xnor (d105, d51, d59);
	buf (d106, d37);
	and (d107, d49, d54);
	buf (d108, d29);
	nor (d109, d47, d77);
	buf (d110, d4);
	nor (d111, d45, d59);
	nand (d112, d64, d75);
	buf (d113, d49);
	nand (d114, d59, d66);
	buf (d115, d69);
	nand (d116, d100, d110);
	not (d117, d81);
	xor (d118, d82, d114);
	buf (d119, d66);
	not (d120, d72);
	assign f1 = d119;
	assign f2 = d117;
	assign f3 = d120;
	assign f4 = d118;
	assign f5 = d118;
	assign f6 = d120;
	assign f7 = d116;
	assign f8 = d119;
	assign f9 = d116;
	assign f10 = d119;
	assign f11 = d119;
	assign f12 = d119;
	assign f13 = d118;
	assign f14 = d119;
	assign f15 = d120;
	assign f16 = d116;
	assign f17 = d120;
	assign f18 = d117;
	assign f19 = d116;
	assign f20 = d119;
endmodule
