module CCGRCG45( x0, x1, x2, x3, f1, f2, f3 );

	input x0, x1, x2, x3;
	output f1, f2, f3;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240;

	not (d1, x1);
	xnor (d2, x3);
	nand (d3, x0, x2);
	nor (d4, x0, x2);
	and (d5, x1, x2);
	nor (d6, x1, x2);
	or (d7, x1, x3);
	xor (d8, x0, x1);
	or (d9, x3);
	nor (d10, x0, x3);
	buf (d11, x2);
	xnor (d12, x0, x1);
	xor (d13, x2, x3);
	xor (d14, x0, x2);
	nand (d15, x1, x2);
	or (d16, x2);
	xnor (d17, x0, x2);
	nor (d18, x2);
	xor (d19, x1, x3);
	and (d20, x0, x1);
	or (d21, x1);
	not (d22, x2);
	nand (d23, x0, x1);
	nand (d24, x1, x2);
	xor (d25, x3);
	nand (d26, x0, x3);
	xnor (d27, x0);
	nor (d28, x0, x1);
	nor (d29, x2, x3);
	buf (d30, x3);
	nor (d31, x3);
	xor (d32, x0);
	or (d33, x2, x3);
	or (d34, x1, x3);
	or (d35, x1, x2);
	xor (d36, x0, x3);
	xor (d37, x2);
	or (d38, x0, x3);
	buf (d39, x0);
	and (d40, x1);
	nand (d41, x2, x3);
	or (d42, x1, x2);
	nand (d43, x0, x1);
	xor (d44, x2, x3);
	and (d45, x1, x2);
	buf (d46, x1);
	nand (d47, x2);
	and (d48, d14, d18);
	or (d49, d13, d41);
	not (d50, d25);
	not (d51, d13);
	nand (d52, d36, d45);
	buf (d53, d42);
	nor (d54, d15, d41);
	nand (d55, d20, d37);
	not (d56, d12);
	and (d57, d9, d20);
	and (d58, d31, d45);
	xor (d59, d17, d30);
	nor (d60, d13, d30);
	and (d61, d30, d42);
	buf (d62, d18);
	and (d63, d9, d45);
	nand (d64, d3, d27);
	nand (d65, d34, d37);
	nand (d66, d61, d65);
	xor (d67, d48, d50);
	xor (d68, d49, d59);
	buf (d69, d41);
	not (d70, d8);
	nor (d71, d56);
	buf (d72, d37);
	buf (d73, d49);
	not (d74, d15);
	xor (d75, d54, d63);
	and (d76, d55, d58);
	or (d77, d51, d65);
	xor (d78, d48, d49);
	and (d79, d49, d57);
	buf (d80, d24);
	nand (d81, d54, d62);
	nor (d82, d52, d55);
	and (d83, d56, d65);
	not (d84, d35);
	nor (d85, d52, d62);
	nor (d86, d58, d65);
	xor (d87, d48, d52);
	and (d88, d54, d61);
	buf (d89, d50);
	and (d90, d56);
	buf (d91, d54);
	and (d92, d59, d63);
	nor (d93, d48, d57);
	nand (d94, d62, d64);
	nand (d95, d56, d60);
	xnor (d96, d60, d63);
	nor (d97, d51, d58);
	or (d98, d50, d58);
	xnor (d99, d61, d65);
	buf (d100, d28);
	and (d101, d48, d64);
	not (d102, d40);
	buf (d103, d1);
	xnor (d104, d60, d64);
	nand (d105, d52, d53);
	nor (d106, d49, d61);
	nor (d107, d52, d57);
	buf (d108, d63);
	not (d109, d46);
	not (d110, d4);
	and (d111, d50, d64);
	buf (d112, d58);
	or (d113, d50, d59);
	not (d114, d27);
	nor (d115, d59, d62);
	nand (d116, d58, d65);
	nand (d117, d58, d61);
	nor (d118, d66, d101);
	not (d119, d34);
	xnor (d120, d71, d84);
	and (d121, d90, d105);
	and (d122, d96, d97);
	nand (d123, d95, d117);
	nand (d124, d68, d117);
	nand (d125, d106);
	and (d126, d78, d98);
	nor (d127, d82, d85);
	and (d128, d96, d101);
	xnor (d129, d105, d109);
	and (d130, d71, d104);
	nand (d131, d94, d116);
	nand (d132, d86, d117);
	not (d133, d5);
	xor (d134, d74, d83);
	or (d135, d85, d100);
	not (d136, d88);
	and (d137, d73, d79);
	and (d138, d84, d104);
	xnor (d139, d69, d108);
	xnor (d140, d82, d83);
	nor (d141, d77, d78);
	nand (d142, d84, d95);
	or (d143, d85, d116);
	and (d144, d75, d102);
	not (d145, d104);
	nor (d146, d72, d114);
	xor (d147, d73, d98);
	and (d148, d105, d116);
	buf (d149, d79);
	buf (d150, d72);
	and (d151, d85, d101);
	nor (d152, d74, d84);
	and (d153, d87, d109);
	nor (d154, d87, d91);
	or (d155, d83, d115);
	nand (d156, d77, d94);
	not (d157, d107);
	nor (d158, d71, d81);
	xor (d159, d93, d100);
	nand (d160, d96, d113);
	nor (d161, d98, d107);
	and (d162, d86, d90);
	xnor (d163, d96, d109);
	not (d164, d81);
	xor (d165, d66, d82);
	and (d166, d99, d101);
	not (d167, d106);
	xnor (d168, d77, d98);
	and (d169, d89, d116);
	xnor (d170, d95, d112);
	xnor (d171, d83, d110);
	or (d172, d67, d90);
	xnor (d173, d111);
	or (d174, d67, d99);
	nor (d175, d105, d107);
	xnor (d176, d86, d89);
	xnor (d177, d101, d104);
	buf (d178, d21);
	not (d179, d48);
	and (d180, d136, d170);
	nor (d181, d165, d170);
	or (d182, d118, d155);
	not (d183, d162);
	nand (d184, d128, d151);
	not (d185, d135);
	or (d186, d145, d163);
	and (d187, d136, d174);
	xnor (d188, d144, d177);
	nor (d189, d118, d157);
	buf (d190, d176);
	xnor (d191, d134, d164);
	buf (d192, d48);
	nand (d193, d137);
	or (d194, d156, d168);
	and (d195, d149, d164);
	xor (d196, d123, d139);
	nand (d197, d147, d162);
	xnor (d198, d131, d153);
	nor (d199, d154, d163);
	xnor (d200, d161, d178);
	and (d201, d135, d151);
	or (d202, d120, d175);
	xnor (d203, d157, d178);
	nand (d204, d134, d165);
	xor (d205, d157, d173);
	and (d206, d147, d172);
	nor (d207, d124, d144);
	nor (d208, d132, d151);
	nor (d209, d167, d168);
	and (d210, d157, d158);
	xor (d211, d125, d164);
	nor (d212, d148, d152);
	nor (d213, d140, d152);
	nand (d214, d136, d162);
	and (d215, d136, d148);
	nor (d216, d157, d158);
	buf (d217, d153);
	nor (d218, d143, d159);
	xor (d219, d133, d157);
	xnor (d220, d137, d157);
	xnor (d221, d172, d174);
	nor (d222, d138, d165);
	nor (d223, d123, d150);
	xnor (d224, d129, d138);
	xor (d225, d141, d173);
	xor (d226, d147, d168);
	or (d227, d148, d169);
	and (d228, d126, d128);
	buf (d229, d139);
	buf (d230, d110);
	and (d231, d122, d157);
	not (d232, d43);
	not (d233, d124);
	nand (d234, d138, d151);
	xor (d235, d132, d163);
	and (d236, d124, d176);
	nor (d237, d152, d174);
	xnor (d238, d130, d142);
	xnor (d239, d152, d173);
	nor (d240, d152, d156);
	assign f1 = d187;
	assign f2 = d229;
	assign f3 = d221;
endmodule
