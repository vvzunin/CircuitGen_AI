module CCGRCG13( x0, x1, f1, f2, f3, f4, f5, f6, f7, f8 );

	input x0, x1;
	output f1, f2, f3, f4, f5, f6, f7, f8;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107;

	not (d1, x1);
	not (d2, x0);
	or (d3, x0, x1);
	nor (d4, x1);
	nand (d5, x0);
	xnor (d6, x0, x1);
	xor (d7, x1);
	and (d8, x1);
	xnor (d9, x0, x1);
	buf (d10, x0);
	xor (d11, x0, x1);
	xnor (d12, x0);
	and (d13, x0, x1);
	or (d14, x0, x1);
	nor (d15, x0, x1);
	and (d16, x0);
	buf (d17, x1);
	xnor (d18, x1);
	nand (d19, x0, x1);
	nor (d20, x0);
	and (d21, x0, x1);
	xor (d22, x0, x1);
	nand (d23, x0, x1);
	nor (d24, x0, x1);
	or (d25, x1);
	xor (d26, x0);
	nand (d27, x1);
	xor (d28, d12, d21);
	xnor (d29, d11, d24);
	xor (d30, d7, d11);
	xnor (d31, d3, d24);
	nand (d32, d14, d20);
	and (d33, d3, d26);
	nand (d34, d6, d12);
	xnor (d35, d22, d26);
	nand (d36, d5, d11);
	xor (d37, d10, d19);
	and (d38, d4, d20);
	not (d39, d18);
	nand (d40, d8, d19);
	xnor (d41, d1, d18);
	buf (d42, d22);
	xor (d43, d16, d25);
	nand (d44, d4, d11);
	xor (d45, d5, d8);
	not (d46, d14);
	not (d47, d8);
	nand (d48, d7, d17);
	or (d49, d6, d24);
	nand (d50, d12, d20);
	or (d51, d4, d14);
	xor (d52, d10, d22);
	nand (d53, d8, d20);
	xor (d54, d27);
	nor (d55, d8, d23);
	xnor (d56, d2, d12);
	not (d57, d17);
	or (d58, d6, d15);
	and (d59, d6, d7);
	not (d60, d7);
	not (d61, d10);
	xor (d62, d10, d11);
	and (d63, d21, d24);
	or (d64, d13, d18);
	and (d65, d6);
	and (d66, d3, d27);
	nor (d67, d25, d26);
	or (d68, d5, d23);
	buf (d69, d26);
	xnor (d70, d1, d25);
	nand (d71, d7, d20);
	and (d72, d1, d8);
	nand (d73, d11, d25);
	and (d74, d3, d23);
	nand (d75, d7, d12);
	xnor (d76, d3, d15);
	xor (d77, d1, d24);
	nand (d78, d7, d25);
	buf (d79, d12);
	buf (d80, d4);
	or (d81, d6, d14);
	or (d82, d3, d21);
	and (d83, d2, d21);
	xnor (d84, d7, d17);
	or (d85, d2, d21);
	xnor (d86, d16, d17);
	not (d87, d27);
	not (d88, d21);
	nor (d89, d11, d21);
	nor (d90, d21, d25);
	buf (d91, d18);
	and (d92, d2, d6);
	nand (d93, d13, d25);
	nand (d94, d15, d23);
	or (d95, d4, d27);
	nor (d96, d23, d24);
	not (d97, d23);
	xor (d98, d18, d19);
	xnor (d99, d15);
	nand (d100, d19, d24);
	nand (d101, d1, d26);
	and (d102, d11, d15);
	nand (d103, d9, d23);
	nand (d104, d4, d14);
	xnor (d105, d12, d27);
	and (d106, d7, d11);
	or (d107, d12, d23);
	assign f1 = d28;
	assign f2 = d66;
	assign f3 = d82;
	assign f4 = d47;
	assign f5 = d39;
	assign f6 = d103;
	assign f7 = d45;
	assign f8 = d102;
endmodule
