module CCGRCG36( x0, x1, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17, f18, f19, f20 );

	input x0, x1;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17, f18, f19, f20;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314, d315, d316, d317, d318, d319, d320, d321, d322, d323, d324, d325, d326, d327, d328, d329, d330, d331, d332, d333, d334, d335, d336, d337, d338, d339, d340, d341, d342, d343, d344, d345, d346, d347, d348, d349, d350, d351, d352, d353, d354, d355, d356, d357, d358, d359, d360, d361, d362, d363, d364, d365, d366, d367, d368, d369, d370, d371, d372, d373, d374, d375, d376, d377, d378, d379, d380, d381, d382, d383, d384, d385, d386, d387, d388, d389, d390, d391, d392, d393, d394, d395, d396, d397, d398, d399, d400, d401, d402, d403, d404, d405, d406, d407, d408, d409, d410, d411, d412, d413, d414, d415, d416, d417, d418, d419, d420, d421, d422, d423, d424, d425, d426, d427, d428, d429, d430, d431, d432, d433, d434, d435, d436, d437, d438, d439, d440, d441, d442, d443, d444, d445, d446, d447, d448, d449, d450, d451, d452, d453, d454, d455, d456, d457, d458, d459, d460, d461, d462, d463, d464, d465, d466, d467, d468, d469, d470, d471, d472, d473, d474, d475, d476, d477, d478, d479, d480, d481, d482, d483, d484, d485, d486, d487, d488, d489, d490, d491, d492, d493, d494, d495, d496, d497, d498, d499, d500, d501, d502, d503, d504, d505, d506, d507, d508, d509, d510, d511, d512, d513, d514, d515, d516, d517, d518, d519, d520, d521, d522, d523, d524, d525, d526, d527, d528, d529, d530, d531, d532, d533, d534, d535, d536, d537, d538, d539, d540, d541, d542, d543, d544, d545, d546, d547, d548, d549, d550, d551, d552, d553, d554, d555, d556, d557, d558, d559, d560, d561, d562, d563, d564, d565, d566, d567, d568, d569, d570, d571, d572, d573, d574, d575, d576, d577, d578, d579, d580, d581, d582, d583, d584, d585, d586, d587, d588;

	or (d1, x0);
	xor (d2, x0);
	not (d3, x0);
	nand (d4, x0, x1);
	xnor (d5, x0);
	buf (d6, x0);
	or (d7, x0, x1);
	and (d8, x0, x1);
	not (d9, x1);
	nand (d10, x0);
	nor (d11, x0);
	xnor (d12, x0, x1);
	nand (d13, x1);
	and (d14, x0);
	xor (d15, x0, x1);
	nor (d16, x1);
	buf (d17, x1);
	nor (d18, x0, x1);
	and (d19, x0, x1);
	xnor (d20, x1);
	or (d21, x1);
	nand (d22, x0, x1);
	xor (d23, x1);
	and (d24, x1);
	xnor (d25, x0, x1);
	nor (d26, x0, x1);
	xor (d27, d6, d11);
	or (d28, d20, d26);
	and (d29, d4, d20);
	or (d30, d2, d3);
	buf (d31, d16);
	or (d32, d11, d25);
	not (d33, d11);
	xnor (d34, d4, d9);
	nor (d35, d21, d24);
	xnor (d36, d5, d21);
	xor (d37, d4, d26);
	nand (d38, d1, d13);
	xnor (d39, d16, d25);
	buf (d40, d7);
	xnor (d41, d2, d6);
	xor (d42, d1, d13);
	not (d43, d17);
	xor (d44, d4, d13);
	xor (d45, d1, d3);
	not (d46, d9);
	nor (d47, d3, d17);
	buf (d48, d25);
	nand (d49, d7, d9);
	buf (d50, d20);
	nand (d51, d16);
	not (d52, d22);
	or (d53, d4, d22);
	xor (d54, d9, d16);
	xor (d55, d7, d15);
	xor (d56, d18, d26);
	xor (d57, d12, d25);
	not (d58, d2);
	nor (d59, d4, d20);
	or (d60, d2, d16);
	nor (d61, d17, d21);
	and (d62, d1, d13);
	nor (d63, d19, d22);
	nor (d64, d8, d24);
	nor (d65, d16, d19);
	xnor (d66, d3, d23);
	and (d67, d2, d26);
	nand (d68, d11, d22);
	or (d69, d8, d9);
	and (d70, d1, d15);
	buf (d71, d8);
	nor (d72, d2, d15);
	not (d73, d10);
	nand (d74, d2, d15);
	not (d75, d8);
	nor (d76, d2, d12);
	buf (d77, d6);
	nand (d78, d14, d24);
	not (d79, d20);
	xor (d80, d4, d19);
	nor (d81, d7, d24);
	not (d82, d14);
	nand (d83, d5, d9);
	and (d84, d4, d14);
	xnor (d85, d11, d21);
	nand (d86, d12);
	nand (d87, d19, d21);
	nand (d88, d7, d12);
	buf (d89, d17);
	nor (d90, d12, d23);
	xor (d91, d20, d25);
	and (d92, d3, d4);
	nor (d93, d12, d19);
	buf (d94, d1);
	nand (d95, d4, d8);
	xnor (d96, d24);
	not (d97, d25);
	nand (d98, d13);
	nand (d99, d9, d17);
	xnor (d100, d9, d22);
	and (d101, d6, d23);
	and (d102, d9, d13);
	xor (d103, d1, d8);
	nor (d104, d17, d23);
	or (d105, d5, d10);
	and (d106, d6, d24);
	xor (d107, d1, d6);
	nand (d108, d22, d23);
	xor (d109, d21, d22);
	and (d110, d6, d18);
	xnor (d111, d15, d24);
	xnor (d112, d9, d18);
	and (d113, d2, d13);
	buf (d114, d13);
	nor (d115, d38, d57);
	nand (d116, d37, d80);
	or (d117, d54, d104);
	or (d118, d54, d104);
	xnor (d119, d86, d101);
	and (d120, d52, d77);
	or (d121, d49, d111);
	and (d122, d39, d41);
	not (d123, d108);
	xor (d124, d84, d114);
	nand (d125, d30, d110);
	or (d126, d68, d75);
	or (d127, d32, d58);
	not (d128, d78);
	nor (d129, d37, d106);
	or (d130, d43, d85);
	nand (d131, d83, d86);
	xnor (d132, d74, d97);
	and (d133, d46, d59);
	and (d134, d110);
	xor (d135, d30, d38);
	nor (d136, d55, d88);
	not (d137, d40);
	xnor (d138, d44, d71);
	nor (d139, d34, d55);
	xnor (d140, d41, d70);
	nand (d141, d39, d104);
	xnor (d142, d60, d87);
	xnor (d143, d77, d94);
	not (d144, d72);
	nand (d145, d34, d103);
	and (d146, d45, d75);
	xnor (d147, d69, d99);
	xnor (d148, d50, d106);
	or (d149, d82, d87);
	xor (d150, d75, d81);
	and (d151, d42, d84);
	and (d152, d51, d95);
	xnor (d153, d45, d103);
	nand (d154, d90, d99);
	nor (d155, d36, d54);
	xor (d156, d47, d99);
	xor (d157, d67, d96);
	or (d158, d38, d73);
	or (d159, d65, d83);
	and (d160, d69, d91);
	or (d161, d52, d57);
	nor (d162, d37, d75);
	and (d163, d93, d101);
	xnor (d164, d85, d108);
	or (d165, d41, d60);
	nand (d166, d47, d107);
	xor (d167, d36, d52);
	nor (d168, d29, d59);
	and (d169, d62, d69);
	buf (d170, d111);
	xnor (d171, d36, d44);
	or (d172, d68, d104);
	nor (d173, d28, d47);
	buf (d174, d135);
	nand (d175, d116, d142);
	buf (d176, d158);
	xor (d177, d136, d159);
	buf (d178, d85);
	xor (d179, d120, d137);
	and (d180, d133, d163);
	nor (d181, d137, d147);
	and (d182, d141, d148);
	buf (d183, d133);
	xor (d184, d146, d156);
	or (d185, d119, d128);
	nand (d186, d149, d172);
	not (d187, d26);
	xor (d188, d117, d160);
	not (d189, d85);
	nor (d190, d152, d153);
	and (d191, d135, d167);
	or (d192, d127, d143);
	nand (d193, d153, d164);
	xor (d194, d158, d169);
	nand (d195, d118, d138);
	not (d196, d106);
	nor (d197, d154, d171);
	xor (d198, d176, d178);
	nand (d199, d179, d188);
	xnor (d200, d175, d194);
	nor (d201, d185, d186);
	xnor (d202, d188, d190);
	nor (d203, d175, d195);
	xnor (d204, d187, d188);
	not (d205, d161);
	or (d206, d176, d181);
	not (d207, d139);
	xor (d208, d176, d195);
	xor (d209, d184, d195);
	nor (d210, d176, d195);
	or (d211, d183, d189);
	nand (d212, d191, d192);
	xor (d213, d183, d187);
	xnor (d214, d174, d197);
	or (d215, d189, d193);
	nor (d216, d175, d176);
	xnor (d217, d178, d190);
	or (d218, d177, d190);
	nor (d219, d181, d191);
	or (d220, d188, d192);
	or (d221, d181, d193);
	xor (d222, d190, d193);
	nor (d223, d195);
	and (d224, d178, d184);
	or (d225, d176, d178);
	or (d226, d184, d187);
	nor (d227, d184, d192);
	not (d228, d23);
	or (d229, d182, d193);
	and (d230, d177, d182);
	nand (d231, d190, d192);
	xnor (d232, d177, d195);
	not (d233, d69);
	not (d234, d46);
	xor (d235, d183);
	nand (d236, d177, d192);
	nor (d237, d186, d189);
	nand (d238, d185, d194);
	xor (d239, d185, d190);
	not (d240, d159);
	not (d241, d175);
	xor (d242, d174, d189);
	nand (d243, d175, d184);
	nand (d244, d176, d191);
	xor (d245, d187, d189);
	buf (d246, d31);
	nor (d247, d183, d194);
	or (d248, d177, d181);
	or (d249, d177, d189);
	buf (d250, d173);
	xor (d251, d186, d193);
	nand (d252, d176, d197);
	nor (d253, d191, d192);
	or (d254, d183, d185);
	xor (d255, d182, d188);
	xor (d256, d174, d184);
	or (d257, d187);
	not (d258, d61);
	nor (d259, d202, d253);
	xor (d260, d237, d238);
	xnor (d261, d253, d256);
	and (d262, d222, d251);
	xor (d263, d235, d236);
	buf (d264, d255);
	xor (d265, d249, d255);
	xnor (d266, d208, d243);
	xor (d267, d199, d239);
	or (d268, d241, d258);
	not (d269, d49);
	or (d270, d219, d240);
	or (d271, d210, d211);
	xor (d272, d202, d240);
	nor (d273, d234, d240);
	xnor (d274, d229, d237);
	buf (d275, d145);
	not (d276, d158);
	xnor (d277, d204, d207);
	or (d278, d201, d257);
	and (d279, d220, d246);
	not (d280, d256);
	nand (d281, d227, d233);
	or (d282, d211, d250);
	nor (d283, d205, d253);
	xnor (d284, d206, d214);
	xnor (d285, d222, d239);
	not (d286, d60);
	nor (d287, d219, d243);
	xnor (d288, d231, d234);
	xnor (d289, d201, d209);
	xor (d290, d198, d220);
	not (d291, d32);
	xnor (d292, d219, d256);
	and (d293, d202, d226);
	buf (d294, d22);
	xnor (d295, d246, d248);
	not (d296, d202);
	nor (d297, d228, d244);
	nand (d298, d200, d227);
	xor (d299, d240, d242);
	nand (d300, d227, d230);
	xor (d301, d210, d240);
	xnor (d302, d225, d251);
	nor (d303, d227, d245);
	nor (d304, d198, d250);
	nand (d305, d215, d226);
	xor (d306, d214, d250);
	xnor (d307, d202, d203);
	buf (d308, d132);
	buf (d309, d121);
	xor (d310, d234, d250);
	or (d311, d235, d244);
	xor (d312, d218, d239);
	or (d313, d205);
	and (d314, d206, d239);
	xnor (d315, d225, d250);
	nand (d316, d218, d220);
	buf (d317, d142);
	nand (d318, d216, d235);
	xor (d319, d212, d254);
	not (d320, d70);
	xnor (d321, d204, d231);
	or (d322, d203, d230);
	nand (d323, d224, d244);
	xnor (d324, d246, d251);
	nand (d325, d205, d247);
	nor (d326, d219, d236);
	or (d327, d249, d258);
	and (d328, d201, d227);
	nand (d329, d253, d255);
	xnor (d330, d244, d251);
	nor (d331, d200, d229);
	nand (d332, d214, d243);
	not (d333, d109);
	or (d334, d206, d223);
	nand (d335, d225, d240);
	buf (d336, d78);
	buf (d337, d62);
	xor (d338, d212, d245);
	or (d339, d216, d249);
	nor (d340, d206, d207);
	xor (d341, d228, d244);
	or (d342, d198, d249);
	xnor (d343, d203, d235);
	xor (d344, d237, d256);
	buf (d345, d149);
	buf (d346, d80);
	and (d347, d238, d243);
	not (d348, d112);
	not (d349, d186);
	nor (d350, d212, d250);
	xor (d351, d255, d258);
	nand (d352, d213, d227);
	nand (d353, d225, d244);
	nand (d354, d263, d309);
	xor (d355, d281, d312);
	and (d356, d336);
	and (d357, d313, d326);
	xnor (d358, d260, d332);
	buf (d359, d213);
	not (d360, d297);
	xor (d361, d303, d350);
	xnor (d362, d292, d294);
	and (d363, d268, d335);
	buf (d364, d146);
	xnor (d365, d259, d270);
	buf (d366, d242);
	xor (d367, d287, d330);
	nand (d368, d340, d342);
	buf (d369, d244);
	nand (d370, d307, d334);
	nor (d371, d263, d281);
	and (d372, d301, d319);
	buf (d373, d353);
	buf (d374, d101);
	not (d375, d250);
	nand (d376, d281, d315);
	nor (d377, d261, d322);
	and (d378, d264, d272);
	buf (d379, d296);
	or (d380, d263, d319);
	not (d381, d88);
	xnor (d382, d268, d351);
	not (d383, d172);
	and (d384, d263, d298);
	xor (d385, d267, d349);
	or (d386, d267, d288);
	nand (d387, d276, d282);
	nand (d388, d259, d328);
	and (d389, d335, d346);
	and (d390, d288, d329);
	not (d391, d248);
	xnor (d392, d296, d315);
	xnor (d393, d286, d320);
	xor (d394, d334, d348);
	and (d395, d264, d316);
	nand (d396, d317, d345);
	nor (d397, d267, d285);
	nor (d398, d285, d349);
	and (d399, d292, d342);
	not (d400, d157);
	nand (d401, d310, d334);
	not (d402, d128);
	nand (d403, d315, d352);
	nor (d404, d324, d343);
	buf (d405, d11);
	nor (d406, d262, d301);
	buf (d407, d307);
	or (d408, d298, d344);
	xnor (d409, d297, d298);
	xor (d410, d293, d296);
	xnor (d411, d301, d324);
	buf (d412, d208);
	or (d413, d292, d343);
	nor (d414, d314, d336);
	buf (d415, d76);
	and (d416, d320, d335);
	or (d417, d275, d311);
	xnor (d418, d305, d334);
	buf (d419, d67);
	not (d420, d211);
	xnor (d421, d288, d313);
	or (d422, d263, d344);
	not (d423, d98);
	and (d424, d275, d306);
	and (d425, d290, d331);
	xor (d426, d325, d331);
	nor (d427, d284, d313);
	not (d428, d253);
	and (d429, d279, d283);
	xnor (d430, d290, d314);
	and (d431, d293, d301);
	nand (d432, d283, d340);
	xnor (d433, d324, d345);
	xor (d434, d288, d336);
	or (d435, d277, d345);
	xor (d436, d292, d300);
	xor (d437, d270, d275);
	xor (d438, d280, d322);
	and (d439, d342, d353);
	buf (d440, d210);
	nand (d441, d296, d350);
	xnor (d442, d264, d280);
	nor (d443, d287, d303);
	not (d444, d113);
	and (d445, d305, d332);
	or (d446, d309, d350);
	buf (d447, d316);
	xor (d448, d312, d332);
	nor (d449, d264, d336);
	xnor (d450, d307, d333);
	or (d451, d269, d318);
	buf (d452, d261);
	xor (d453, d395, d400);
	buf (d454, d216);
	or (d455, d395, d399);
	xor (d456, d389, d425);
	buf (d457, d385);
	not (d458, d412);
	xnor (d459, d426, d449);
	buf (d460, d407);
	and (d461, d363, d418);
	or (d462, d410, d436);
	buf (d463, d390);
	not (d464, d93);
	or (d465, d367, d440);
	and (d466, d365, d387);
	and (d467, d444, d450);
	xor (d468, d365, d376);
	nor (d469, d415, d443);
	not (d470, d147);
	xnor (d471, d405, d437);
	and (d472, d402, d436);
	xor (d473, d397, d405);
	nand (d474, d390, d419);
	buf (d475, d379);
	xnor (d476, d406, d413);
	not (d477, d372);
	not (d478, d429);
	xnor (d479, d399, d440);
	xor (d480, d364, d376);
	nand (d481, d379, d392);
	and (d482, d405, d413);
	nand (d483, d363, d371);
	and (d484, d358, d424);
	xor (d485, d414, d428);
	nor (d486, d373, d446);
	xor (d487, d401, d450);
	xor (d488, d376, d386);
	xor (d489, d398, d451);
	xor (d490, d355, d429);
	xnor (d491, d416, d426);
	xnor (d492, d395, d404);
	or (d493, d405, d438);
	xor (d494, d361, d392);
	xnor (d495, d358, d440);
	not (d496, d384);
	xnor (d497, d359, d415);
	or (d498, d443, d446);
	nor (d499, d369, d380);
	not (d500, d5);
	nor (d501, d405, d416);
	xor (d502, d394, d447);
	buf (d503, d23);
	not (d504, d255);
	xor (d505, d395, d410);
	nand (d506, d380, d385);
	and (d507, d459, d466);
	buf (d508, d300);
	not (d509, d337);
	nand (d510, d454, d485);
	xor (d511, d480, d494);
	or (d512, d455, d489);
	nand (d513, d470, d492);
	nand (d514, d460, d474);
	nor (d515, d475, d480);
	xor (d516, d480, d488);
	nand (d517, d482, d484);
	buf (d518, d322);
	xor (d519, d490, d493);
	buf (d520, d372);
	xor (d521, d489, d498);
	xor (d522, d454, d490);
	nand (d523, d456, d484);
	not (d524, d19);
	not (d525, d35);
	nand (d526, d457, d500);
	xor (d527, d463, d464);
	and (d528, d470, d479);
	nand (d529, d468, d474);
	nor (d530, d480, d505);
	not (d531, d154);
	nand (d532, d466, d498);
	nand (d533, d458, d469);
	xor (d534, d472, d473);
	nand (d535, d485, d493);
	nand (d536, d473, d476);
	xor (d537, d486, d504);
	or (d538, d457, d498);
	xnor (d539, d453, d492);
	and (d540, d468, d488);
	and (d541, d480, d482);
	nor (d542, d453, d472);
	xor (d543, d489, d496);
	and (d544, d495, d497);
	nor (d545, d474, d477);
	nand (d546, d455, d496);
	nor (d547, d458, d475);
	buf (d548, d402);
	not (d549, d185);
	xor (d550, d464, d502);
	xor (d551, d473, d475);
	buf (d552, d271);
	and (d553, d488, d495);
	buf (d554, d168);
	nor (d555, d478, d496);
	xnor (d556, d484, d499);
	nand (d557, d479, d491);
	nor (d558, d490, d494);
	nand (d559, d504, d505);
	nor (d560, d484, d489);
	and (d561, d482, d496);
	xor (d562, d459, d506);
	and (d563, d460, d481);
	or (d564, d461, d496);
	xor (d565, d453, d465);
	buf (d566, d114);
	not (d567, d181);
	buf (d568, d479);
	nand (d569, d461, d506);
	xnor (d570, d481, d487);
	xnor (d571, d461, d505);
	nand (d572, d482, d501);
	or (d573, d463, d503);
	buf (d574, d219);
	xor (d575, d454, d505);
	nor (d576, d478, d505);
	not (d577, d210);
	xnor (d578, d485, d489);
	nor (d579, d457, d483);
	buf (d580, d10);
	and (d581, d478, d493);
	nor (d582, d489, d493);
	nor (d583, d456, d471);
	and (d584, d460, d465);
	xnor (d585, d473, d502);
	nor (d586, d493, d505);
	or (d587, d476, d477);
	nand (d588, d455, d484);
	assign f1 = d521;
	assign f2 = d526;
	assign f3 = d564;
	assign f4 = d540;
	assign f5 = d584;
	assign f6 = d541;
	assign f7 = d536;
	assign f8 = d584;
	assign f9 = d513;
	assign f10 = d509;
	assign f11 = d559;
	assign f12 = d572;
	assign f13 = d569;
	assign f14 = d552;
	assign f15 = d545;
	assign f16 = d552;
	assign f17 = d536;
	assign f18 = d525;
	assign f19 = d514;
	assign f20 = d509;
endmodule
