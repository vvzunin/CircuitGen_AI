module CCGRCG104( x0, x1, x2, x3, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16 );

	input x0, x1, x2, x3;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314, d315, d316, d317, d318, d319, d320, d321, d322, d323, d324, d325, d326;

	xor (d1, x0, x1);
	buf (d2, x3);
	not (d3, x3);
	nor (d4, x2, x3);
	or (d5, x1, x3);
	and (d6, x0, x2);
	buf (d7, x1);
	and (d8, x0, x1);
	xnor (d9, x0, x3);
	xnor (d10, x2);
	and (d11, x0, x3);
	or (d12, x0, x2);
	xnor (d13, x0);
	buf (d14, x2);
	xnor (d15, d1, d4);
	not (d16, d12);
	nor (d17, d6, d9);
	not (d18, d5);
	nand (d19, d4, d6);
	xnor (d20, d4, d12);
	nand (d21, d3, d6);
	and (d22, d7, d12);
	xor (d23, d1, d14);
	xnor (d24, d3, d14);
	xnor (d25, d4, d5);
	buf (d26, d4);
	nand (d27, d12, d14);
	xor (d28, d1, d7);
	and (d29, d3, d4);
	or (d30, d3, d14);
	nand (d31, d3, d11);
	nor (d32, d2, d10);
	nor (d33, d10, d13);
	and (d34, d13, d14);
	buf (d35, d10);
	not (d36, d14);
	buf (d37, d8);
	not (d38, x1);
	xnor (d39, d9, d13);
	or (d40, d8, d11);
	buf (d41, d11);
	xor (d42, d2, d4);
	not (d43, d7);
	not (d44, x0);
	nand (d45, d1, d6);
	and (d46, d9, d14);
	and (d47, d11, d14);
	and (d48, d2, d5);
	and (d49, d8, d12);
	xor (d50, d6);
	xor (d51, d3);
	xor (d52, d2, d11);
	buf (d53, d3);
	not (d54, d1);
	nand (d55, d10, d12);
	nor (d56, d1, d11);
	or (d57, d5, d11);
	and (d58, d2, d10);
	buf (d59, d9);
	and (d60, d11, d14);
	or (d61, d4, d14);
	and (d62, d3, d5);
	xor (d63, d5, d14);
	and (d64, d2, d12);
	xnor (d65, d2, d6);
	and (d66, d9, d10);
	or (d67, d3, d13);
	nand (d68, d1, d2);
	xnor (d69, d35, d65);
	not (d70, d24);
	buf (d71, d35);
	nand (d72, d17, d40);
	and (d73, d38, d49);
	xor (d74, d16, d45);
	xnor (d75, d44, d62);
	xnor (d76, d22, d59);
	buf (d77, d41);
	xnor (d78, d31, d63);
	xor (d79, d38, d40);
	or (d80, d33, d62);
	xnor (d81, d25, d48);
	or (d82, d18, d35);
	or (d83, d28, d39);
	xnor (d84, d46, d49);
	not (d85, d34);
	and (d86, d22, d54);
	or (d87, d35, d48);
	or (d88, d40);
	or (d89, d20, d40);
	xor (d90, d18, d59);
	xnor (d91, d24, d58);
	nor (d92, d41, d42);
	xnor (d93, d24, d64);
	and (d94, d48, d52);
	xnor (d95, d15, d16);
	and (d96, d17, d35);
	nor (d97, d17, d26);
	xnor (d98, d36, d43);
	or (d99, d36, d53);
	buf (d100, d39);
	nor (d101, d42, d59);
	buf (d102, d19);
	nand (d103, d30, d62);
	or (d104, d51, d59);
	xnor (d105, d46, d51);
	xnor (d106, d46, d58);
	xor (d107, d23, d48);
	or (d108, d55);
	nor (d109, d52, d56);
	xnor (d110, d47, d59);
	nor (d111, d25, d67);
	not (d112, d65);
	nor (d113, d17, d67);
	nand (d114, d15, d34);
	nand (d115, d48, d63);
	not (d116, x2);
	nor (d117, d20, d36);
	or (d118, d31, d34);
	xnor (d119, d66, d68);
	buf (d120, d34);
	xnor (d121, d22, d52);
	and (d122, d44, d64);
	nand (d123, d39, d63);
	xor (d124, d39, d53);
	nor (d125, d15, d50);
	or (d126, d29, d32);
	xnor (d127, d44, d53);
	xor (d128, d48, d60);
	nor (d129, d19, d25);
	nor (d130, d49, d59);
	xor (d131, d21, d24);
	and (d132, d40, d57);
	nand (d133, d40, d68);
	or (d134, d25, d52);
	xnor (d135, d30, d37);
	nand (d136, d19, d68);
	nor (d137, d31, d33);
	or (d138, d50, d68);
	nand (d139, d33, d41);
	xnor (d140, d43, d63);
	xor (d141, d32, d62);
	not (d142, d38);
	xor (d143, d48, d50);
	or (d144, d28, d62);
	and (d145, d29, d68);
	nor (d146, d49);
	or (d147, d27, d65);
	and (d148, d40, d62);
	nand (d149, d18, d30);
	buf (d150, d7);
	xor (d151, d23, d60);
	not (d152, d6);
	and (d153, d44, d60);
	nand (d154, d49, d65);
	or (d155, d37, d53);
	and (d156, d30, d36);
	not (d157, d8);
	and (d158, d27, d65);
	xor (d159, d70, d83);
	not (d160, d91);
	and (d161, d94, d115);
	xor (d162, d145, d149);
	nand (d163, d83, d147);
	or (d164, d124, d132);
	xnor (d165, d119, d154);
	buf (d166, d57);
	buf (d167, d70);
	or (d168, d152, d154);
	xnor (d169, d102, d134);
	and (d170, d75, d82);
	or (d171, d77, d147);
	or (d172, d116, d138);
	or (d173, d115, d127);
	not (d174, d41);
	or (d175, d112, d150);
	or (d176, d84, d114);
	xor (d177, d81, d158);
	xor (d178, d70, d80);
	buf (d179, d133);
	or (d180, d73, d131);
	buf (d181, d152);
	buf (d182, d149);
	xnor (d183, d99, d110);
	buf (d184, d12);
	nand (d185, d101, d139);
	buf (d186, d150);
	not (d187, d135);
	nand (d188, d81, d122);
	or (d189, d69, d127);
	xnor (d190, d118, d146);
	or (d191, d130, d140);
	and (d192, d88, d95);
	nand (d193, d92, d149);
	xnor (d194, d127, d142);
	or (d195, d95, d151);
	xor (d196, d108, d137);
	not (d197, d28);
	xnor (d198, d100, d127);
	nor (d199, d122, d155);
	not (d200, d70);
	and (d201, d83, d127);
	xnor (d202, d104, d110);
	xor (d203, d117, d118);
	and (d204, d74, d107);
	xnor (d205, d91, d119);
	not (d206, d51);
	nand (d207, d74, d155);
	xnor (d208, d146, d147);
	nor (d209, d101, d120);
	or (d210, d82, d149);
	buf (d211, d104);
	nor (d212, d120, d140);
	not (d213, d50);
	nor (d214, d183, d204);
	or (d215, d170, d195);
	buf (d216, d203);
	xor (d217, d176, d189);
	nand (d218, d174, d211);
	not (d219, d73);
	and (d220, d181, d200);
	nor (d221, d165, d173);
	nor (d222, d166, d179);
	or (d223, d187, d209);
	nand (d224, d175, d182);
	nor (d225, d159, d188);
	not (d226, d152);
	or (d227, d164, d200);
	and (d228, d178, d190);
	and (d229, d180, d184);
	nand (d230, d185, d201);
	xnor (d231, d162, d185);
	and (d232, d163, d167);
	nand (d233, d191, d202);
	xnor (d234, d161, d204);
	and (d235, d165, d203);
	xnor (d236, d188, d198);
	or (d237, d172, d186);
	nand (d238, d166, d192);
	xnor (d239, d180, d207);
	nor (d240, d167, d195);
	nand (d241, d204, d210);
	or (d242, d179, d213);
	nor (d243, d191, d194);
	xor (d244, d205, d211);
	xor (d245, d197, d208);
	not (d246, d121);
	and (d247, d172, d186);
	buf (d248, d182);
	buf (d249, d15);
	or (d250, d161, d204);
	nand (d251, d161, d210);
	xor (d252, d179, d203);
	xnor (d253, d224);
	nor (d254, d214, d224);
	xor (d255, d248, d250);
	buf (d256, d186);
	xor (d257, d240, d250);
	and (d258, d235, d241);
	xnor (d259, d214, d250);
	nor (d260, d239, d246);
	nand (d261, d219, d220);
	xor (d262, d214, d240);
	xnor (d263, d231, d246);
	buf (d264, d160);
	xnor (d265, d232);
	nand (d266, d232, d248);
	xor (d267, d237, d241);
	and (d268, d225, d244);
	xor (d269, d223, d249);
	buf (d270, d67);
	nor (d271, d226, d232);
	xnor (d272, d245, d248);
	or (d273, d219, d249);
	or (d274, d220, d247);
	xnor (d275, d225, d243);
	xnor (d276, d231, d237);
	nor (d277, d216, d234);
	nand (d278, d218, d235);
	and (d279, d225, d250);
	xnor (d280, d223, d241);
	nand (d281, d226, d242);
	xor (d282, d220, d237);
	buf (d283, d137);
	xnor (d284, d217, d225);
	or (d285, d249, d250);
	xnor (d286, d236, d243);
	and (d287, d237, d244);
	nand (d288, d222, d239);
	and (d289, d216, d240);
	or (d290, d215, d225);
	nand (d291, d228, d242);
	xnor (d292, d233, d251);
	xor (d293, d235, d246);
	xnor (d294, d220, d232);
	buf (d295, d227);
	not (d296, d105);
	nor (d297, d226, d245);
	not (d298, d110);
	or (d299, d214, d235);
	xnor (d300, d216, d247);
	xnor (d301, d224, d228);
	nor (d302, d235, d242);
	buf (d303, d217);
	xor (d304, d229, d233);
	not (d305, d78);
	xnor (d306, d229, d232);
	xor (d307, d243, d252);
	or (d308, d224, d242);
	or (d309, d235, d250);
	xnor (d310, d237, d242);
	not (d311, d36);
	xnor (d312, d221, d243);
	xor (d313, d235, d239);
	buf (d314, d231);
	and (d315, d231, d238);
	or (d316, d222, d244);
	and (d317, d228, d233);
	xnor (d318, d231, d249);
	not (d319, d184);
	and (d320, d230, d241);
	or (d321, d223, d250);
	xnor (d322, d229, d252);
	buf (d323, d183);
	nor (d324, d217, d225);
	nor (d325, d231, d242);
	xnor (d326, d227, d248);
	assign f1 = d269;
	assign f2 = d325;
	assign f3 = d320;
	assign f4 = d262;
	assign f5 = d321;
	assign f6 = d279;
	assign f7 = d258;
	assign f8 = d260;
	assign f9 = d265;
	assign f10 = d258;
	assign f11 = d278;
	assign f12 = d289;
	assign f13 = d295;
	assign f14 = d324;
	assign f15 = d277;
	assign f16 = d263;
endmodule
