module CCGRCG67( x0, x1, x2, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16 );

	input x0, x1, x2;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38;

	and (d1, x0, x2);
	nand (d2, x0);
	xor (d3, x1, x2);
	xor (d4, x2);
	or (d5, x0, x2);
	and (d6, x2);
	not (d7, x0);
	nor (d8, x1, x2);
	xor (d9, x0, x1);
	xnor (d10, x0);
	not (d11, x1);
	xor (d12, x0, x2);
	buf (d13, x2);
	or (d14, x2);
	xnor (d15, x0, x2);
	nand (d16, x2);
	nor (d17, x0, x1);
	nand (d18, x1, x2);
	nor (d19, x2);
	not (d20, x2);
	xor (d21, x1, x2);
	and (d22, x1);
	nand (d23, x0, x2);
	xor (d24, x1);
	and (d25, x0);
	xnor (d26, x1, x2);
	xor (d27, x0, x2);
	and (d28, x1, x2);
	nor (d29, x1, x2);
	xnor (d30, x1, x2);
	and (d31, x0, x1);
	or (d32, x0, x1);
	buf (d33, x1);
	xor (d34, x0, x1);
	or (d35, x1, x2);
	xnor (d36, x0, x1);
	and (d37, x1, x2);
	or (d38, x0, x1);
	assign f1 = d20;
	assign f2 = d1;
	assign f3 = d1;
	assign f4 = d4;
	assign f5 = d37;
	assign f6 = d27;
	assign f7 = d3;
	assign f8 = d5;
	assign f9 = d26;
	assign f10 = d18;
	assign f11 = d3;
	assign f12 = d29;
	assign f13 = d27;
	assign f14 = d23;
	assign f15 = d18;
	assign f16 = d5;
endmodule
