module CCGRCG16( x0, x1, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10 );

	input x0, x1;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200;

	nand (d1, x1);
	or (d2, x0, x1);
	xnor (d3, x0, x1);
	not (d4, x1);
	and (d5, x0);
	buf (d6, x0);
	and (d7, x0, x1);
	buf (d8, x1);
	nor (d9, x0, x1);
	nand (d10, x0, x1);
	xor (d11, x0);
	xnor (d12, x1);
	nor (d13, x1);
	or (d14, x0, x1);
	not (d15, x0);
	nand (d16, x0);
	and (d17, x0, x1);
	or (d18, x1);
	xor (d19, x1);
	nor (d20, x0);
	nor (d21, x0, x1);
	and (d22, x1);
	xor (d23, x0, x1);
	or (d24, x0);
	xnor (d25, x0, x1);
	nand (d26, x0, x1);
	xnor (d27, x0);
	xnor (d28, d23, d25);
	nor (d29, d3, d8);
	nand (d30, d10, d11);
	or (d31, d5, d17);
	or (d32, d5, d25);
	buf (d33, d11);
	or (d34, d9, d15);
	xor (d35, d14, d18);
	xor (d36, d1, d5);
	or (d37, d2, d10);
	nor (d38, d19, d21);
	nor (d39, d1, d5);
	not (d40, d25);
	and (d41, d9, d26);
	not (d42, d3);
	xnor (d43, d2, d16);
	nor (d44, d4, d16);
	xor (d45, d13, d16);
	xnor (d46, d6, d7);
	or (d47, d5, d9);
	and (d48, d4, d9);
	nor (d49, d4, d27);
	and (d50, d15, d18);
	xnor (d51, d2, d13);
	and (d52, d16, d25);
	nand (d53, d1, d7);
	not (d54, d11);
	nand (d55, d5, d13);
	nand (d56, d25, d27);
	nor (d57, d47, d55);
	and (d58, d35, d46);
	and (d59, d51, d56);
	buf (d60, d15);
	and (d61, d56);
	nand (d62, d35, d56);
	xor (d63, d37, d43);
	nand (d64, d29, d33);
	nor (d65, d39, d49);
	buf (d66, d21);
	nor (d67, d46, d56);
	or (d68, d32, d55);
	buf (d69, d45);
	xor (d70, d32, d34);
	xor (d71, d32, d56);
	nand (d72, d29, d35);
	nor (d73, d32, d45);
	nand (d74, d38, d53);
	or (d75, d49, d50);
	nand (d76, d44, d54);
	nand (d77, d36, d52);
	and (d78, d40, d46);
	xnor (d79, d57, d77);
	xnor (d80, d76, d78);
	not (d81, d68);
	xnor (d82, d68, d69);
	buf (d83, d26);
	or (d84, d64, d78);
	xor (d85, d71, d77);
	or (d86, d74, d75);
	not (d87, d50);
	xor (d88, d66, d72);
	nor (d89, d66, d70);
	xor (d90, d59, d60);
	nand (d91, d61, d70);
	buf (d92, d64);
	or (d93, d63, d68);
	or (d94, d58, d64);
	or (d95, d63, d70);
	xor (d96, d67, d74);
	nor (d97, d67, d69);
	nand (d98, d65, d77);
	nor (d99, d59, d77);
	xor (d100, d67, d76);
	nand (d101, d57, d58);
	nor (d102, d67, d71);
	nor (d103, d61, d66);
	nand (d104, d62, d72);
	nor (d105, d65, d76);
	nor (d106, d72, d74);
	xor (d107, d61, d68);
	buf (d108, d6);
	buf (d109, d50);
	not (d110, d26);
	nor (d111, d64, d66);
	xnor (d112, d57, d77);
	xor (d113, d69, d71);
	xor (d114, d64, d75);
	not (d115, d65);
	buf (d116, d46);
	xnor (d117, d64, d68);
	nand (d118, d93, d105);
	or (d119, d101, d110);
	nand (d120, d82, d97);
	nor (d121, d99, d107);
	xnor (d122, d82, d93);
	and (d123, d88, d102);
	nor (d124, d107, d112);
	or (d125, d90, d95);
	not (d126, d66);
	and (d127, d98, d104);
	buf (d128, d36);
	xor (d129, d92, d107);
	and (d130, d86, d101);
	and (d131, d97, d101);
	buf (d132, d62);
	buf (d133, d28);
	xor (d134, d90, d93);
	xnor (d135, d97, d99);
	nand (d136, d81, d116);
	nor (d137, d85, d104);
	or (d138, d97, d116);
	buf (d139, d52);
	or (d140, d86, d98);
	and (d141, d83, d100);
	or (d142, d87, d92);
	xor (d143, d124, d129);
	not (d144, d40);
	not (d145, d113);
	or (d146, d119, d127);
	buf (d147, d114);
	xor (d148, d125, d139);
	and (d149, d133, d135);
	not (d150, d86);
	nor (d151, d130, d137);
	and (d152, d125, d142);
	xor (d153, d132, d133);
	nor (d154, d136, d140);
	and (d155, d125, d142);
	xnor (d156, d121, d136);
	and (d157, d122, d141);
	buf (d158, d83);
	nor (d159, d135, d137);
	xor (d160, d123, d131);
	nor (d161, d130, d136);
	nor (d162, d130, d138);
	and (d163, d137, d141);
	nor (d164, d128, d134);
	or (d165, d133, d137);
	not (d166, d135);
	or (d167, d121, d130);
	or (d168, d127, d129);
	nand (d169, d125, d137);
	xor (d170, d127, d131);
	or (d171, d124, d125);
	and (d172, d120, d123);
	xor (d173, d130, d133);
	and (d174, d131, d141);
	or (d175, d121, d136);
	xnor (d176, d124, d141);
	or (d177, d120, d132);
	buf (d178, d125);
	or (d179, d130, d138);
	not (d180, d38);
	and (d181, d119, d123);
	buf (d182, d105);
	nor (d183, d131, d135);
	or (d184, d118, d133);
	or (d185, d118, d125);
	nor (d186, d120, d139);
	nand (d187, d131, d139);
	xor (d188, d122, d140);
	buf (d189, d110);
	nand (d190, d121);
	not (d191, d111);
	nand (d192, d119, d121);
	not (d193, d121);
	not (d194, d55);
	nand (d195, d121, d131);
	or (d196, d118, d122);
	not (d197, d17);
	or (d198, d122, d142);
	nand (d199, d125, d128);
	buf (d200, d106);
	assign f1 = d156;
	assign f2 = d156;
	assign f3 = d179;
	assign f4 = d183;
	assign f5 = d191;
	assign f6 = d188;
	assign f7 = d197;
	assign f8 = d197;
	assign f9 = d189;
	assign f10 = d193;
endmodule
