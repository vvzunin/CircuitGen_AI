module CCGRCG40( x0, x1, x2, x3, f1 );

	input x0, x1, x2, x3;
	output f1;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74;

	buf (d1, x3);
	xnor (d2, x3);
	or (d3, x1, x3);
	nand (d4, x2, x3);
	nand (d5, x0, x1);
	and (d6, x0);
	nor (d7, x2, x3);
	nand (d8, x2, x3);
	buf (d9, x2);
	or (d10, x0, x3);
	buf (d11, x0);
	xnor (d12, x0, x3);
	and (d13, x2, x3);
	and (d14, x2, x3);
	and (d15, x1, x2);
	not (d16, x1);
	xnor (d17, x0);
	not (d18, x0);
	or (d19, x2, x3);
	not (d20, x2);
	xnor (d21, x0, x2);
	nand (d22, x0, x2);
	xor (d23, x2, x3);
	or (d24, x0, x2);
	or (d25, x2, x3);
	or (d26, x3);
	nor (d27, x1, x2);
	and (d28, x0, x2);
	xor (d29, x1, x2);
	buf (d30, x1);
	or (d31, x0, x1);
	or (d32, x0, x1);
	xnor (d33, x1, x2);
	xnor (d34, x2, x3);
	and (d35, d7, d24);
	buf (d36, d27);
	buf (d37, d33);
	xnor (d38, d10, d22);
	xor (d39, d11, d19);
	xor (d40, d15, d29);
	nand (d41, d3, d11);
	not (d42, d15);
	buf (d43, d10);
	nand (d44, d6, d16);
	nand (d45, d13);
	buf (d46, d17);
	buf (d47, d15);
	xnor (d48, d28, d33);
	not (d49, d9);
	not (d50, d30);
	not (d51, d1);
	or (d52, d5, d19);
	nor (d53, d3, d9);
	nand (d54, d19, d33);
	and (d55, d2, d8);
	not (d56, d4);
	and (d57, d4, d21);
	nand (d58, d7, d33);
	xnor (d59, d7, d30);
	nand (d60, d21, d28);
	nand (d61, d16, d32);
	xnor (d62, d6, d10);
	nand (d63, d6, d21);
	nand (d64, d15, d32);
	nand (d65, d9);
	not (d66, d20);
	nand (d67, d33, d34);
	nor (d68, d22, d31);
	nor (d69, d21, d30);
	xor (d70, d11, d14);
	nand (d71, d14, d20);
	and (d72, d29, d33);
	xor (d73, d22, d27);
	nor (d74, d26);
	assign f1 = d64;
endmodule
