module CCGRCG35( x0, x1, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17, f18, f19 );

	input x0, x1;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17, f18, f19;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314, d315, d316, d317, d318, d319, d320, d321, d322, d323, d324, d325, d326, d327, d328, d329, d330, d331, d332, d333, d334, d335, d336, d337, d338, d339, d340, d341, d342, d343, d344, d345, d346, d347, d348, d349, d350, d351, d352, d353, d354, d355, d356, d357, d358, d359, d360, d361, d362, d363, d364, d365, d366, d367, d368, d369, d370, d371, d372, d373, d374, d375, d376, d377, d378, d379, d380, d381, d382, d383, d384, d385, d386, d387, d388, d389, d390, d391, d392, d393, d394, d395, d396, d397, d398, d399, d400, d401, d402, d403, d404, d405, d406, d407, d408, d409, d410, d411, d412, d413, d414, d415, d416, d417, d418, d419, d420, d421, d422, d423, d424;

	nand (d1, x0);
	and (d2, x0, x1);
	xnor (d3, x1);
	nand (d4, x1);
	or (d5, d1, d3);
	and (d6, d1, d3);
	buf (d7, d3);
	and (d8, d3, d4);
	nand (d9, d1, d2);
	nor (d10, d3);
	buf (d11, x1);
	or (d12, d4);
	xnor (d13, d3);
	nor (d14, d1);
	xor (d15, d1, d2);
	or (d16, d2, d3);
	nand (d17, d3, d4);
	or (d18, d1, d3);
	xnor (d19, d1, d4);
	xnor (d20, d2);
	or (d21, d2, d4);
	nor (d22, d2, d4);
	or (d23, d1, d4);
	nand (d24, d2);
	and (d25, d2, d4);
	and (d26, d1, d4);
	not (d27, d3);
	not (d28, x1);
	xor (d29, d2, d4);
	xnor (d30, d1, d2);
	xor (d31, d2, d4);
	nor (d32, d3, d4);
	nand (d33, d1, d4);
	xor (d34, d1, d3);
	xnor (d35, d1, d2);
	or (d36, d1, d2);
	or (d37, d3, d4);
	nor (d38, d1, d4);
	nor (d39, d1, d2);
	nand (d40, d2, d3);
	nand (d41, d1, d3);
	xor (d42, d3, d4);
	nand (d43, d3);
	xnor (d44, d1, d3);
	nor (d45, d1, d4);
	or (d46, d2);
	not (d47, d1);
	or (d48, d2, d4);
	or (d49, d1, d2);
	and (d50, d1, d3);
	buf (d51, d1);
	xnor (d52, d3, d4);
	not (d53, d4);
	xor (d54, d1);
	nand (d55, d2, d4);
	or (d56, d1, d4);
	not (d57, x0);
	not (d58, d2);
	xnor (d59, d2, d3);
	xor (d60, d3, d4);
	buf (d61, d2);
	buf (d62, d29);
	nand (d63, d26, d27);
	not (d64, d55);
	nor (d65, d21, d34);
	nor (d66, d18, d20);
	and (d67, d11, d58);
	nand (d68, d22, d43);
	and (d69, d66);
	not (d70, d30);
	xor (d71, d67);
	xor (d72, d65, d66);
	and (d73, d62, d65);
	not (d74, d61);
	xnor (d75, d64, d67);
	not (d76, d59);
	xor (d77, d64, d65);
	xor (d78, d63, d65);
	xor (d79, d62, d66);
	or (d80, d66, d68);
	nor (d81, d62, d65);
	buf (d82, d60);
	xor (d83, d64, d68);
	xor (d84, d66);
	not (d85, d15);
	xor (d86, d63, d67);
	or (d87, d66, d68);
	not (d88, d60);
	and (d89, d65);
	or (d90, d66, d67);
	not (d91, d35);
	xor (d92, d63, d67);
	or (d93, d67, d68);
	xor (d94, d64, d66);
	and (d95, d62, d67);
	buf (d96, d20);
	or (d97, d62, d65);
	nor (d98, d62, d63);
	buf (d99, d14);
	xnor (d100, d62, d67);
	not (d101, d33);
	xnor (d102, d62, d68);
	and (d103, d66, d67);
	or (d104, d62, d68);
	or (d105, d62);
	xor (d106, d68);
	nand (d107, d63, d68);
	or (d108, d65, d68);
	xnor (d109, d66);
	nand (d110, d67);
	nor (d111, d63);
	xor (d112, d64, d65);
	nor (d113, d62, d66);
	not (d114, d13);
	buf (d115, d25);
	xnor (d116, d63, d66);
	xnor (d117, d66, d68);
	not (d118, d65);
	nor (d119, d64, d65);
	or (d120, d62, d63);
	not (d121, d41);
	nand (d122, d64, d67);
	nand (d123, d63, d64);
	or (d124, d64, d65);
	and (d125, d65, d67);
	xnor (d126, d64, d65);
	and (d127, d64);
	buf (d128, d38);
	or (d129, d65, d66);
	and (d130, d67);
	xnor (d131, d66, d67);
	not (d132, d25);
	xor (d133, d62, d65);
	xnor (d134, d65, d66);
	or (d135, d62, d64);
	nor (d136, d65, d68);
	xnor (d137, d65);
	xnor (d138, d64, d68);
	buf (d139, d37);
	nand (d140, d67, d68);
	nand (d141, d63, d67);
	xor (d142, d66, d67);
	not (d143, d19);
	nor (d144, d62, d65);
	nor (d145, d64, d68);
	buf (d146, d16);
	nor (d147, d66);
	and (d148, d115, d141);
	nor (d149, d105, d140);
	xor (d150, d78, d126);
	nand (d151, d77, d125);
	buf (d152, d81);
	not (d153, d49);
	nand (d154, d91, d106);
	xor (d155, d69, d128);
	or (d156, d70, d122);
	nand (d157, d100, d110);
	or (d158, d86, d94);
	xor (d159, d75, d125);
	nor (d160, d76, d99);
	xor (d161, d126, d127);
	not (d162, d136);
	nand (d163, d76, d129);
	nor (d164, d100, d130);
	or (d165, d72, d142);
	nand (d166, d83, d107);
	nor (d167, d103, d106);
	nand (d168, d82, d135);
	xor (d169, d71, d76);
	nor (d170, d97, d145);
	or (d171, d97, d117);
	xor (d172, d111, d130);
	buf (d173, d56);
	xnor (d174, d94, d141);
	not (d175, d16);
	or (d176, d107, d128);
	xor (d177, d77, d84);
	not (d178, d132);
	nand (d179, d95, d100);
	or (d180, d106, d137);
	nand (d181, d79, d120);
	nand (d182, d132, d136);
	nor (d183, d98, d113);
	nand (d184, d72, d126);
	not (d185, d106);
	nand (d186, d72);
	not (d187, d115);
	nor (d188, d85, d110);
	and (d189, d133, d137);
	and (d190, d96, d119);
	xnor (d191, d85, d136);
	and (d192, d83, d108);
	xnor (d193, d93, d99);
	nor (d194, d116, d129);
	xnor (d195, d74, d113);
	xnor (d196, d104, d132);
	or (d197, d78, d122);
	xor (d198, d101, d102);
	nand (d199, d81, d110);
	nand (d200, d94, d134);
	nor (d201, d90, d134);
	not (d202, d74);
	xnor (d203, d140, d142);
	nand (d204, d119, d126);
	or (d205, d93, d121);
	xor (d206, d108, d113);
	not (d207, d31);
	or (d208, d105, d133);
	buf (d209, d102);
	and (d210, d120, d127);
	nand (d211, d133, d147);
	not (d212, d40);
	xnor (d213, d97, d108);
	and (d214, d88, d99);
	or (d215, d78, d131);
	nor (d216, d87, d126);
	nor (d217, d79, d129);
	xor (d218, d101, d120);
	and (d219, d139, d146);
	or (d220, d77, d113);
	not (d221, d119);
	buf (d222, d104);
	and (d223, d106, d118);
	xor (d224, d99, d145);
	nand (d225, d72, d106);
	not (d226, d116);
	buf (d227, d8);
	nor (d228, d185, d190);
	or (d229, d176, d192);
	and (d230, d154, d197);
	xor (d231, d149, d215);
	nor (d232, d174, d196);
	xor (d233, d195, d213);
	buf (d234, d153);
	or (d235, d175, d207);
	xnor (d236, d174, d197);
	nand (d237, d191, d225);
	and (d238, d170, d196);
	xnor (d239, d184, d223);
	or (d240, d157, d184);
	buf (d241, d100);
	nand (d242, d179, d182);
	xnor (d243, d157, d167);
	xor (d244, d199, d205);
	xnor (d245, d168, d197);
	nand (d246, d174, d216);
	not (d247, d166);
	and (d248, d177, d192);
	buf (d249, d202);
	xor (d250, d210, d216);
	or (d251, d213, d216);
	xor (d252, d148, d163);
	not (d253, d6);
	buf (d254, d147);
	or (d255, d172, d212);
	nand (d256, d191, d207);
	not (d257, d184);
	nor (d258, d235, d237);
	xor (d259, d251, d255);
	not (d260, d205);
	and (d261, d234, d235);
	and (d262, d248, d251);
	xnor (d263, d233, d235);
	xor (d264, d241, d251);
	xor (d265, d229, d239);
	and (d266, d252, d255);
	or (d267, d231, d242);
	nand (d268, d238, d239);
	or (d269, d233, d243);
	nand (d270, d239, d245);
	xnor (d271, d234, d244);
	nand (d272, d250, d251);
	and (d273, d231, d241);
	not (d274, d255);
	nor (d275, d229, d252);
	and (d276, d261, d265);
	nand (d277, d257, d273);
	and (d278, d257, d270);
	not (d279, d248);
	or (d280, d258, d271);
	and (d281, d265, d267);
	xor (d282, d257, d264);
	nor (d283, d260, d268);
	or (d284, d257, d263);
	xnor (d285, d266, d267);
	or (d286, d257, d273);
	nand (d287, d265, d269);
	xnor (d288, d258, d269);
	nor (d289, d260, d264);
	nand (d290, d259, d261);
	not (d291, d66);
	and (d292, d257, d267);
	and (d293, d258, d270);
	or (d294, d266, d268);
	xnor (d295, d260, d269);
	nand (d296, d274, d275);
	nor (d297, d257, d265);
	or (d298, d266, d267);
	or (d299, d262, d265);
	xnor (d300, d258, d268);
	or (d301, d257, d263);
	xnor (d302, d266, d273);
	and (d303, d276, d285);
	nor (d304, d292, d302);
	not (d305, d45);
	nor (d306, d283, d297);
	not (d307, d201);
	and (d308, d280, d292);
	and (d309, d279, d288);
	and (d310, d292, d300);
	nor (d311, d276, d281);
	nor (d312, d292, d293);
	or (d313, d293, d302);
	nand (d314, d282, d302);
	nand (d315, d291, d302);
	xor (d316, d295, d298);
	or (d317, d283, d293);
	nor (d318, d291, d296);
	nor (d319, d279, d287);
	or (d320, d280, d291);
	and (d321, d291, d302);
	nand (d322, d282, d291);
	and (d323, d277, d289);
	not (d324, d244);
	nand (d325, d290, d294);
	or (d326, d298, d299);
	and (d327, d295, d301);
	not (d328, d8);
	and (d329, d277, d302);
	and (d330, d286, d299);
	nand (d331, d290, d300);
	not (d332, d71);
	nand (d333, d281, d294);
	xor (d334, d285, d296);
	or (d335, d279, d281);
	nor (d336, d291, d300);
	nor (d337, d278, d287);
	nor (d338, d282, d301);
	or (d339, d279, d293);
	or (d340, d278, d298);
	xnor (d341, d278, d298);
	xnor (d342, d279);
	or (d343, d286, d300);
	and (d344, d296, d302);
	not (d345, d123);
	or (d346, d294, d300);
	buf (d347, d118);
	and (d348, d277, d292);
	xor (d349, d319, d326);
	not (d350, d177);
	not (d351, d77);
	and (d352, d327, d339);
	or (d353, d334, d346);
	and (d354, d307, d319);
	nor (d355, d332, d334);
	nand (d356, d315, d333);
	not (d357, d29);
	or (d358, d335, d340);
	or (d359, d324, d333);
	xor (d360, d333, d346);
	xor (d361, d317, d337);
	and (d362, d308, d312);
	buf (d363, d70);
	buf (d364, d26);
	nor (d365, d306, d346);
	or (d366, d318, d330);
	nand (d367, d311, d314);
	buf (d368, d319);
	xor (d369, d308, d309);
	nand (d370, d308, d343);
	xor (d371, d320, d335);
	nand (d372, d319, d331);
	nor (d373, d328, d338);
	buf (d374, d19);
	xor (d375, d311, d328);
	and (d376, d328, d336);
	buf (d377, d257);
	xnor (d378, d330, d344);
	nand (d379, d313, d321);
	nor (d380, d316, d325);
	xnor (d381, d322, d340);
	or (d382, d310, d337);
	nand (d383, d326, d331);
	or (d384, d317, d347);
	xor (d385, d330, d346);
	not (d386, d197);
	and (d387, d311, d325);
	not (d388, d161);
	nand (d389, d303, d311);
	or (d390, d316, d331);
	nand (d391, d313, d341);
	or (d392, d304, d338);
	and (d393, d337, d341);
	or (d394, d303, d318);
	or (d395, d342, d345);
	buf (d396, d21);
	not (d397, d252);
	nor (d398, d306, d333);
	nor (d399, d331, d337);
	nand (d400, d329, d341);
	xnor (d401, d309, d330);
	not (d402, d52);
	or (d403, d312, d340);
	and (d404, d319, d340);
	nor (d405, d308, d330);
	xnor (d406, d313, d348);
	nand (d407, d318, d323);
	nor (d408, d330, d336);
	buf (d409, d291);
	xor (d410, d308, d335);
	nor (d411, d303, d322);
	not (d412, d254);
	or (d413, d315, d319);
	buf (d414, d231);
	xor (d415, d315, d331);
	or (d416, d305, d314);
	not (d417, d282);
	buf (d418, d234);
	xnor (d419, d312, d341);
	nor (d420, d314, d348);
	or (d421, d318, d331);
	xor (d422, d318, d347);
	and (d423, d319, d345);
	not (d424, d300);
	assign f1 = d408;
	assign f2 = d376;
	assign f3 = d363;
	assign f4 = d375;
	assign f5 = d417;
	assign f6 = d374;
	assign f7 = d384;
	assign f8 = d359;
	assign f9 = d409;
	assign f10 = d357;
	assign f11 = d380;
	assign f12 = d366;
	assign f13 = d421;
	assign f14 = d349;
	assign f15 = d371;
	assign f16 = d386;
	assign f17 = d423;
	assign f18 = d382;
	assign f19 = d349;
endmodule
