module CCGRCG20( x0, x1, x2, f1 );

	input x0, x1, x2;
	output f1;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59;

	xor (d1, x1, x2);
	xnor (d2, x0);
	nand (d3, x0, x1);
	xnor (d4, x1, x2);
	xnor (d5, x0, x1);
	buf (d6, x1);
	buf (d7, x2);
	or (d8, x1);
	nor (d9, x0, x1);
	nor (d10, x0, x2);
	xor (d11, x0, x2);
	not (d12, x0);
	and (d13, x0, x1);
	not (d14, x2);
	xor (d15, x0, x2);
	nor (d16, x1);
	or (d17, x0, x1);
	xnor (d18, x2);
	xor (d19, x0);
	xor (d20, x0, x1);
	buf (d21, x0);
	nand (d22, x1, x2);
	nor (d23, x0, x1);
	nand (d24, x2);
	xnor (d25, x0, x2);
	nand (d26, x0, x1);
	or (d27, x1, x2);
	and (d28, x1, x2);
	or (d29, x0, x1);
	nor (d30, x1, x2);
	nand (d31, x0, x2);
	nand (d32, x1, x2);
	xnor (d33, x0, x1);
	or (d34, x1, x2);
	and (d35, x0, x2);
	or (d36, x0);
	xor (d37, x1);
	or (d38, x0, x2);
	nor (d39, x0, x2);
	nor (d40, x2);
	nor (d41, x0);
	not (d42, x1);
	xor (d43, x0, x1);
	not (d44, d28);
	nand (d45, d18, d21);
	nor (d46, d2, d13);
	xor (d47, d10, d24);
	nor (d48, d26, d27);
	or (d49, d30);
	nor (d50, d29, d43);
	nor (d51, d7, d32);
	and (d52, d8, d37);
	xnor (d53, d7, d40);
	xor (d54, d1, d17);
	xor (d55, d4, d25);
	buf (d56, d42);
	buf (d57, d33);
	xnor (d58, d8, d20);
	xor (d59, d3, d38);
	assign f1 = d49;
endmodule
