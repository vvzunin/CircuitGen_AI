module CCGRCG133( x0, x1, x2, x3, x4, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11 );

	input x0, x1, x2, x3, x4;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314, d315, d316, d317, d318, d319, d320, d321, d322, d323, d324, d325, d326, d327, d328, d329, d330, d331, d332, d333, d334, d335, d336, d337, d338, d339, d340, d341, d342, d343, d344, d345, d346, d347, d348, d349, d350, d351, d352, d353, d354, d355, d356, d357, d358, d359, d360, d361, d362, d363, d364, d365, d366, d367, d368, d369, d370;

	buf (d1, x3);
	not (d2, x1);
	buf (d3, x2);
	xnor (d4, x1, x3);
	or (d5, x0, x1);
	xnor (d6, x0, x4);
	not (d7, x2);
	xnor (d8, x1, x4);
	not (d9, x3);
	nor (d10, x1, x4);
	nor (d11, x2, x4);
	xnor (d12, x4);
	buf (d13, x1);
	buf (d14, x0);
	or (d15, x2, x3);
	not (d16, x4);
	xor (d17, x3, x4);
	xnor (d18, x1, x3);
	or (d19, x3);
	or (d20, x0, x4);
	xor (d21, x0, x4);
	or (d22, x0, x3);
	and (d23, x0, x3);
	buf (d24, x4);
	nor (d25, x1, x3);
	or (d26, x0, x2);
	xnor (d27, x1, x4);
	or (d28, x4);
	or (d29, x0, x3);
	nor (d30, x3, x4);
	nand (d31, x0, x2);
	or (d32, x0, x2);
	xnor (d33, x0, x4);
	or (d34, x2, x3);
	or (d35, x1, x2);
	nor (d36, x1, x2);
	nor (d37, x0, x4);
	nor (d38, x1, x2);
	nor (d39, x1);
	not (d40, x0);
	xor (d41, x1, x2);
	and (d42, x1, x3);
	nand (d43, x2, x4);
	and (d44, x1, x4);
	buf (d45, d37);
	not (d46, d40);
	not (d47, d15);
	nand (d48, d4, d14);
	nor (d49, d15, d42);
	or (d50, d29, d40);
	or (d51, d25, d29);
	nor (d52, d19, d36);
	xor (d53, d26, d37);
	nor (d54, d10, d19);
	and (d55, d3, d9);
	and (d56, d3, d24);
	xor (d57, d22, d38);
	xor (d58, d17, d42);
	or (d59, d6, d8);
	xor (d60, d14, d37);
	buf (d61, d8);
	and (d62, d21, d32);
	nor (d63, d9, d24);
	buf (d64, d7);
	or (d65, d49, d50);
	and (d66, d45, d46);
	not (d67, d53);
	xor (d68, d56, d61);
	nor (d69, d45, d61);
	nor (d70, d51, d54);
	nand (d71, d57, d61);
	xor (d72, d52, d56);
	buf (d73, d59);
	not (d74, d45);
	xnor (d75, d45, d59);
	xnor (d76, d45, d48);
	xnor (d77, d58, d59);
	buf (d78, d52);
	and (d79, d46, d51);
	or (d80, d46, d47);
	xor (d81, d48, d56);
	and (d82, d51, d55);
	and (d83, d47, d52);
	buf (d84, d29);
	nand (d85, d51, d52);
	xnor (d86, d58);
	or (d87, d61);
	buf (d88, d54);
	not (d89, d8);
	nor (d90, d61, d62);
	buf (d91, d19);
	nor (d92, d54, d58);
	buf (d93, d27);
	nor (d94, d46, d59);
	xnor (d95, d50, d59);
	xor (d96, d50, d56);
	not (d97, d5);
	or (d98, d45, d53);
	or (d99, d48, d58);
	or (d100, d50);
	xor (d101, d46, d50);
	nand (d102, d55, d63);
	nor (d103, d50, d54);
	xor (d104, d46);
	buf (d105, d56);
	xor (d106, d48, d52);
	nor (d107, d48, d58);
	xor (d108, d46, d62);
	xnor (d109, d51, d60);
	nand (d110, d57, d59);
	xnor (d111, d57, d61);
	nor (d112, d49);
	xnor (d113, d55, d61);
	or (d114, d52, d55);
	not (d115, d12);
	nor (d116, d61, d63);
	xnor (d117, d55, d56);
	xor (d118, d45, d61);
	nor (d119, d50, d51);
	not (d120, d10);
	xnor (d121, d49, d56);
	not (d122, d2);
	nor (d123, d48, d52);
	nand (d124, d61, d62);
	nand (d125, d56, d58);
	and (d126, d45, d63);
	nor (d127, d45, d57);
	nand (d128, d59, d61);
	nand (d129, d59, d60);
	xnor (d130, d45, d59);
	xnor (d131, d56, d62);
	xnor (d132, d47, d56);
	xnor (d133, d51, d55);
	not (d134, d22);
	or (d135, d61, d62);
	or (d136, d47, d51);
	buf (d137, d42);
	nor (d138, d46, d53);
	nor (d139, d48, d54);
	not (d140, d46);
	nand (d141, d47, d57);
	nand (d142, d47, d50);
	xor (d143, d57, d60);
	not (d144, d38);
	or (d145, d97, d109);
	xor (d146, d69, d130);
	or (d147, d103, d140);
	xor (d148, d89, d130);
	nand (d149, d112, d115);
	and (d150, d66, d111);
	and (d151, d85, d126);
	not (d152, d130);
	nand (d153, d67, d115);
	or (d154, d68, d74);
	nand (d155, d86, d103);
	or (d156, d90, d119);
	not (d157, d72);
	buf (d158, d118);
	and (d159, d113, d127);
	xor (d160, d72, d101);
	xnor (d161, d122, d128);
	nand (d162, d80, d126);
	nor (d163, d81, d143);
	buf (d164, d121);
	buf (d165, d109);
	nor (d166, d136, d137);
	and (d167, d68, d129);
	xnor (d168, d107, d140);
	nor (d169, d91, d127);
	xnor (d170, d94, d116);
	xor (d171, d120, d123);
	or (d172, d94, d106);
	not (d173, d108);
	buf (d174, d139);
	nand (d175, d103, d142);
	nor (d176, d84, d101);
	nor (d177, d82, d106);
	xor (d178, d79, d93);
	xor (d179, d68, d106);
	xnor (d180, d91, d135);
	and (d181, d106, d142);
	buf (d182, d141);
	xor (d183, d76, d101);
	buf (d184, d47);
	nor (d185, d86, d134);
	or (d186, d115, d122);
	nor (d187, d71, d72);
	xor (d188, d97, d121);
	xnor (d189, d69, d97);
	or (d190, d91, d111);
	nor (d191, d65, d116);
	nand (d192, d67, d134);
	not (d193, d144);
	buf (d194, d5);
	nand (d195, d80, d123);
	not (d196, d98);
	and (d197, d82, d130);
	xor (d198, d78, d135);
	nand (d199, d106, d127);
	nand (d200, d75, d88);
	xor (d201, d77, d111);
	buf (d202, d25);
	xnor (d203, d95, d120);
	and (d204, d115, d132);
	or (d205, d86, d111);
	nand (d206, d104, d140);
	xor (d207, d109, d141);
	nand (d208, d99, d111);
	buf (d209, d112);
	nand (d210, d113, d117);
	or (d211, d134, d139);
	xnor (d212, d92, d97);
	or (d213, d82, d93);
	not (d214, d126);
	or (d215, d84, d120);
	xnor (d216, d96, d128);
	nor (d217, d123, d126);
	xor (d218, d105, d122);
	and (d219, d123, d135);
	buf (d220, d105);
	xor (d221, d67, d102);
	and (d222, d101, d108);
	or (d223, d138, d144);
	xor (d224, d74, d135);
	not (d225, d54);
	nor (d226, d66, d128);
	and (d227, d69, d124);
	xor (d228, d93, d119);
	and (d229, d113, d142);
	or (d230, d67, d73);
	buf (d231, d38);
	xnor (d232, d88, d97);
	not (d233, d41);
	or (d234, d109, d130);
	xnor (d235, d81, d143);
	xor (d236, d139, d142);
	xnor (d237, d64, d65);
	not (d238, d120);
	xor (d239, d162, d223);
	nand (d240, d151, d161);
	xor (d241, d164, d177);
	nor (d242, d153, d237);
	and (d243, d149);
	xor (d244, d147, d183);
	not (d245, d57);
	nand (d246, d205, d212);
	buf (d247, d11);
	and (d248, d149, d191);
	nand (d249, d182, d228);
	xor (d250, d173, d189);
	buf (d251, d89);
	and (d252, d220, d222);
	xor (d253, d183, d185);
	and (d254, d154, d156);
	xor (d255, d158, d208);
	and (d256, d151, d216);
	buf (d257, d236);
	nor (d258, d175, d229);
	or (d259, d180, d225);
	nand (d260, d172, d174);
	xor (d261, d146, d173);
	nand (d262, d164, d170);
	nor (d263, d145, d216);
	or (d264, d169, d226);
	xor (d265, d226);
	and (d266, d180, d230);
	xnor (d267, d167, d184);
	xnor (d268, d164, d175);
	xor (d269, d170, d224);
	xnor (d270, d240, d246);
	nor (d271, d239, d260);
	or (d272, d256, d263);
	nand (d273, d241, d258);
	not (d274, d185);
	xor (d275, d246, d251);
	xor (d276, d243, d252);
	buf (d277, d111);
	or (d278, d239, d259);
	nand (d279, d243, d258);
	xnor (d280, d244, d252);
	not (d281, d150);
	xnor (d282, d252, d257);
	buf (d283, d67);
	and (d284, d246, d264);
	and (d285, d272, d284);
	and (d286, d271, d282);
	buf (d287, d93);
	nand (d288, d274, d280);
	or (d289, d275, d276);
	nor (d290, d275, d278);
	and (d291, d275, d276);
	xor (d292, d282, d283);
	nor (d293, d273, d277);
	or (d294, d273, d274);
	not (d295, d100);
	xor (d296, d270, d277);
	xor (d297, d280, d283);
	nand (d298, d278, d284);
	or (d299, d284);
	buf (d300, d120);
	nand (d301, d272, d283);
	or (d302, d270, d274);
	nor (d303, d271, d279);
	xor (d304, d279, d281);
	xnor (d305, d278, d283);
	nand (d306, d280, d282);
	xnor (d307, d271, d274);
	xnor (d308, d277, d284);
	and (d309, d278);
	buf (d310, d106);
	and (d311, d272);
	nor (d312, d271, d274);
	xor (d313, d272, d282);
	and (d314, d284);
	not (d315, d279);
	not (d316, d66);
	nor (d317, d272, d273);
	not (d318, d37);
	buf (d319, d280);
	not (d320, d68);
	and (d321, d271, d279);
	xor (d322, d280);
	or (d323, d273, d277);
	and (d324, d277, d280);
	xor (d325, d270, d278);
	not (d326, d114);
	buf (d327, d281);
	xnor (d328, d275, d276);
	or (d329, d279, d284);
	nand (d330, d274, d284);
	xnor (d331, d272, d280);
	xnor (d332, d281, d283);
	buf (d333, d74);
	buf (d334, d176);
	xnor (d335, d279, d283);
	nand (d336, d275, d281);
	xor (d337, d270, d273);
	nand (d338, d270, d282);
	nand (d339, d274);
	or (d340, d274, d277);
	and (d341, d274, d280);
	and (d342, d273, d274);
	xor (d343, d277, d279);
	xor (d344, d274, d279);
	xnor (d345, d275, d278);
	xnor (d346, d290, d329);
	xnor (d347, d301, d320);
	xnor (d348, d302, d307);
	nor (d349, d290, d321);
	xnor (d350, d291, d307);
	buf (d351, d276);
	nor (d352, d296, d302);
	and (d353, d311, d328);
	nand (d354, d294, d307);
	and (d355, d349, d351);
	nor (d356, d348, d354);
	not (d357, d18);
	or (d358, d346, d349);
	xnor (d359, d348);
	xor (d360, d346, d353);
	nor (d361, d347, d351);
	nor (d362, d349, d350);
	xor (d363, d350);
	nand (d364, d346, d354);
	not (d365, d186);
	or (d366, d346, d354);
	xnor (d367, d348, d352);
	xor (d368, d346, d347);
	or (d369, d352, d354);
	xnor (d370, d346, d353);
	assign f1 = d360;
	assign f2 = d364;
	assign f3 = d363;
	assign f4 = d363;
	assign f5 = d368;
	assign f6 = d357;
	assign f7 = d359;
	assign f8 = d367;
	assign f9 = d356;
	assign f10 = d361;
	assign f11 = d357;
endmodule
