module CCGRCG99( x0, x1, x2, x3, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13 );

	input x0, x1, x2, x3;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311;

	or (d1, x0);
	not (d2, x1);
	or (d3, x0, x1);
	xnor (d4, x0, x3);
	xor (d5, x2, x3);
	and (d6, x3);
	xor (d7, x2, x3);
	nand (d8, x2, x3);
	and (d9, x0, x2);
	buf (d10, x2);
	not (d11, x0);
	or (d12, x2, x3);
	or (d13, x2);
	xor (d14, x0, x1);
	and (d15, x2);
	buf (d16, x3);
	nand (d17, x0, x2);
	buf (d18, x0);
	xnor (d19, x1, x3);
	buf (d20, x1);
	not (d21, x3);
	or (d22, x1, x2);
	xnor (d23, x1);
	nand (d24, x3);
	or (d25, x0, x3);
	or (d26, x0, x2);
	xnor (d27, x0, x3);
	nand (d28, x0, x3);
	xnor (d29, x3);
	xnor (d30, x0, x1);
	and (d31, x0);
	nand (d32, x0, x1);
	xor (d33, x0, x3);
	not (d34, x2);
	nor (d35, x0, x3);
	xor (d36, x0);
	buf (d37, d32);
	nor (d38, d20, d24);
	and (d39, d23, d35);
	xor (d40, d7, d12);
	not (d41, d31);
	nor (d42, d11, d34);
	xor (d43, d28, d33);
	xnor (d44, d9, d14);
	buf (d45, d18);
	not (d46, d34);
	nand (d47, d4, d15);
	and (d48, d17, d18);
	nand (d49, d30, d35);
	xnor (d50, d5, d6);
	and (d51, d3, d18);
	not (d52, d3);
	nand (d53, d10, d15);
	or (d54, d7, d30);
	xnor (d55, d15, d35);
	xnor (d56, d14, d33);
	xnor (d57, d2, d33);
	not (d58, d19);
	or (d59, d34, d36);
	not (d60, d23);
	or (d61, d14, d21);
	nand (d62, d10, d18);
	xnor (d63, d16, d34);
	nor (d64, d19, d23);
	nor (d65, d5, d28);
	xnor (d66, d20, d24);
	nand (d67, d20, d28);
	nand (d68, d19, d28);
	and (d69, d23, d30);
	or (d70, d6, d17);
	xnor (d71, d5, d27);
	and (d72, d12, d28);
	xor (d73, d14, d22);
	nand (d74, d4, d28);
	xnor (d75, d19, d28);
	nor (d76, d18, d36);
	nand (d77, d21, d23);
	not (d78, d6);
	or (d79, d5, d28);
	nor (d80, d17, d35);
	and (d81, d11, d32);
	xnor (d82, d28, d31);
	xor (d83, d13, d24);
	or (d84, d21, d26);
	nor (d85, d14, d27);
	xor (d86, d4, d10);
	xor (d87, d4, d14);
	nand (d88, d24, d25);
	or (d89, d26, d28);
	and (d90, d15, d26);
	not (d91, d27);
	buf (d92, d35);
	or (d93, d20, d21);
	nand (d94, d29, d30);
	xnor (d95, d5, d10);
	xor (d96, d22, d34);
	nand (d97, d26, d31);
	xor (d98, d18, d19);
	and (d99, d2, d4);
	nand (d100, d26, d32);
	not (d101, d21);
	not (d102, d33);
	and (d103, d15, d23);
	or (d104, d20, d24);
	nor (d105, d6, d27);
	xor (d106, d34, d35);
	nand (d107, d2, d10);
	nor (d108, d29, d36);
	and (d109, d9, d14);
	xnor (d110, d35, d36);
	nand (d111, d11, d15);
	nand (d112, d1, d23);
	xor (d113, d25, d31);
	xnor (d114, d19, d24);
	nor (d115, d4, d11);
	not (d116, d15);
	nand (d117, d3, d15);
	nand (d118, d1, d13);
	xnor (d119, d12, d26);
	or (d120, d32, d34);
	and (d121, d23, d31);
	nand (d122, d9, d36);
	or (d123, d17, d35);
	and (d124, d24, d28);
	or (d125, d14, d31);
	xnor (d126, d62, d69);
	or (d127, d53, d90);
	not (d128, d26);
	nor (d129, d89, d125);
	xor (d130, d48, d97);
	or (d131, d50, d122);
	and (d132, d63, d113);
	buf (d133, d5);
	nand (d134, d39, d102);
	buf (d135, d81);
	buf (d136, d116);
	nor (d137, d44, d79);
	buf (d138, d121);
	or (d139, d100, d112);
	or (d140, d62, d101);
	nor (d141, d59, d63);
	not (d142, d107);
	nor (d143, d53, d123);
	xnor (d144, d61, d63);
	xnor (d145, d37, d121);
	not (d146, d20);
	and (d147, d80, d121);
	or (d148, d72, d96);
	and (d149, d56, d124);
	xor (d150, d55, d103);
	not (d151, d73);
	and (d152, d112, d125);
	or (d153, d89, d110);
	nor (d154, d67, d87);
	and (d155, d38, d97);
	nand (d156, d73, d109);
	xnor (d157, d66, d87);
	xor (d158, d79, d107);
	nand (d159, d82, d118);
	or (d160, d63, d84);
	nor (d161, d82, d119);
	xor (d162, d65, d68);
	nand (d163, d48, d94);
	or (d164, d44, d95);
	nor (d165, d86, d105);
	and (d166, d52, d112);
	and (d167, d56, d58);
	xnor (d168, d55, d80);
	or (d169, d63, d122);
	xnor (d170, d39, d123);
	xor (d171, d46, d63);
	or (d172, d45, d69);
	nor (d173, d42, d50);
	or (d174, d65, d107);
	or (d175, d81, d112);
	not (d176, d18);
	nor (d177, d84, d114);
	xnor (d178, d64, d122);
	xnor (d179, d94, d116);
	nor (d180, d55, d60);
	buf (d181, d113);
	nand (d182, d106, d116);
	buf (d183, d42);
	xor (d184, d111, d120);
	not (d185, d77);
	xnor (d186, d96, d105);
	xor (d187, d61, d125);
	and (d188, d51, d54);
	xnor (d189, d102, d109);
	nor (d190, d57, d114);
	nand (d191, d49, d58);
	and (d192, d101, d108);
	nor (d193, d126, d178);
	buf (d194, d58);
	and (d195, d151, d188);
	not (d196, d53);
	xor (d197, d172, d186);
	xnor (d198, d128, d170);
	not (d199, d97);
	xor (d200, d132, d138);
	or (d201, d142, d187);
	xnor (d202, d169, d192);
	xor (d203, d178, d181);
	nand (d204, d189, d192);
	or (d205, d128, d134);
	nand (d206, d144, d189);
	nor (d207, d146, d174);
	nand (d208, d137, d143);
	nand (d209, d141, d191);
	not (d210, d140);
	or (d211, d178, d183);
	xnor (d212, d144, d175);
	nor (d213, d130);
	nand (d214, d132, d161);
	not (d215, d86);
	nand (d216, d153, d159);
	nor (d217, d130, d169);
	nand (d218, d135, d157);
	and (d219, d149, d180);
	not (d220, d158);
	buf (d221, d48);
	and (d222, d168);
	xor (d223, d144, d161);
	nand (d224, d175, d192);
	xnor (d225, d167, d173);
	buf (d226, d162);
	buf (d227, d141);
	buf (d228, d161);
	or (d229, d141, d191);
	buf (d230, d124);
	and (d231, d171, d178);
	xnor (d232, d128, d133);
	nand (d233, d129, d159);
	xnor (d234, d146, d187);
	or (d235, d140, d190);
	xnor (d236, d130, d169);
	not (d237, d89);
	and (d238, d135, d153);
	not (d239, d172);
	nor (d240, d203, d238);
	not (d241, d188);
	or (d242, d207, d234);
	and (d243, d215, d233);
	xor (d244, d205, d222);
	or (d245, d199, d237);
	or (d246, d193, d220);
	xor (d247, d199, d221);
	and (d248, d227, d229);
	xnor (d249, d200, d222);
	not (d250, d2);
	and (d251, d200, d235);
	nand (d252, d215, d232);
	xnor (d253, d201, d222);
	xnor (d254, d197, d212);
	nor (d255, d226, d228);
	nor (d256, d195, d203);
	buf (d257, d190);
	and (d258, d212, d221);
	or (d259, d204, d215);
	nand (d260, d208, d218);
	xor (d261, d194, d204);
	xnor (d262, d231, d232);
	not (d263, d95);
	and (d264, d209, d210);
	nor (d265, d193, d227);
	xor (d266, d202, d214);
	or (d267, d226, d229);
	or (d268, d195);
	not (d269, d139);
	xnor (d270, d200, d228);
	or (d271, d196, d227);
	xnor (d272, d211, d237);
	or (d273, d201, d206);
	nand (d274, d199, d222);
	xor (d275, d199, d208);
	or (d276, d205, d237);
	not (d277, d126);
	xor (d278, d205, d238);
	xnor (d279, d219, d226);
	xnor (d280, d229, d231);
	and (d281, d230, d235);
	and (d282, d205, d206);
	xnor (d283, d194, d234);
	xor (d284, d193, d204);
	xor (d285, d212, d214);
	nand (d286, d197, d226);
	and (d287, d209, d211);
	xor (d288, d195, d236);
	not (d289, d106);
	xor (d290, d199, d214);
	nand (d291, d197, d236);
	or (d292, d204, d208);
	or (d293, d197, d227);
	buf (d294, d148);
	or (d295, d206, d223);
	or (d296, d198, d232);
	nor (d297, d213, d221);
	nor (d298, d193, d235);
	xnor (d299, d205, d221);
	and (d300, d196, d217);
	buf (d301, d80);
	not (d302, d178);
	not (d303, d63);
	nor (d304, d211, d227);
	or (d305, d214, d226);
	nand (d306, d217, d235);
	xnor (d307, d205, d213);
	xnor (d308, d199, d205);
	nor (d309, d214, d219);
	buf (d310, d70);
	xor (d311, d226, d237);
	assign f1 = d269;
	assign f2 = d240;
	assign f3 = d294;
	assign f4 = d239;
	assign f5 = d279;
	assign f6 = d256;
	assign f7 = d308;
	assign f8 = d242;
	assign f9 = d270;
	assign f10 = d255;
	assign f11 = d304;
	assign f12 = d259;
	assign f13 = d295;
endmodule
