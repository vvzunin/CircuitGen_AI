module CCGRCG61( x0, x1, x2, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13 );

	input x0, x1, x2;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45;

	nand (d1, x1, x2);
	xnor (d2, x0, x2);
	not (d3, x2);
	nor (d4, x0, x1);
	or (d5, x0, x2);
	nor (d6, x0, x2);
	nand (d7, x0, x2);
	or (d8, x1);
	xnor (d9, x1, x2);
	buf (d10, x0);
	nand (d11, x0, x1);
	buf (d12, x2);
	and (d13, x1, x2);
	xor (d14, x0, x1);
	xor (d15, x1);
	xor (d16, x0, x1);
	nand (d17, x0, x2);
	xnor (d18, x2);
	or (d19, x0, x1);
	xnor (d20, x1, x2);
	xnor (d21, x0, x1);
	not (d22, x0);
	or (d23, x1, x2);
	buf (d24, x1);
	nor (d25, x0);
	nand (d26, x0, x1);
	nor (d27, x1, x2);
	not (d28, x1);
	xor (d29, x1, x2);
	xnor (d30, x0);
	nor (d31, x0, x1);
	and (d32, x2);
	and (d33, x0, x2);
	xor (d34, x0, x2);
	and (d35, x0);
	xnor (d36, x0, x1);
	and (d37, x1);
	and (d38, x1, x2);
	nor (d39, x2);
	nor (d40, x1, x2);
	nor (d41, x1);
	nand (d42, x2);
	xor (d43, d33, d35);
	xor (d44, d1, d5);
	xnor (d45, d2);
	assign f1 = d45;
	assign f2 = d45;
	assign f3 = d45;
	assign f4 = d43;
	assign f5 = d45;
	assign f6 = d45;
	assign f7 = d43;
	assign f8 = d45;
	assign f9 = d44;
	assign f10 = d45;
	assign f11 = d44;
	assign f12 = d45;
	assign f13 = d43;
endmodule
