module CCGRCG77( x0, x1, x2, x3, f1, f2 );

	input x0, x1, x2, x3;
	output f1, f2;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307;

	xor (d1, x0, x1);
	xnor (d2, x0, x2);
	nor (d3, x1, x3);
	or (d4, x0);
	and (d5, x1, x3);
	nor (d6, x2, x3);
	or (d7, x3);
	xor (d8, x2, x3);
	xnor (d9, x0);
	xnor (d10, x1, x3);
	and (d11, x2);
	xor (d12, x0, x2);
	not (d13, x3);
	nor (d14, x2);
	xnor (d15, x0, x3);
	not (d16, x0);
	nand (d17, x1);
	and (d18, x0, x3);
	buf (d19, x1);
	nand (d20, x0);
	xor (d21, x1);
	and (d22, x0, x2);
	not (d23, x2);
	xnor (d24, x1, x2);
	or (d25, x1);
	or (d26, x2, x3);
	not (d27, x1);
	nand (d28, x0, x2);
	nor (d29, x1, x2);
	and (d30, x3);
	xnor (d31, x0, x3);
	or (d32, x1, x2);
	nor (d33, x0, x1);
	nand (d34, x1, x3);
	buf (d35, x2);
	or (d36, x1, x3);
	or (d37, x0, x2);
	and (d38, x1, x2);
	nor (d39, d26, d38);
	nor (d40, d6, d36);
	buf (d41, d11);
	xor (d42, d11, d23);
	buf (d43, d22);
	xor (d44, d19, d38);
	xor (d45, d7, d20);
	not (d46, d28);
	nand (d47, d1, d8);
	not (d48, d6);
	buf (d49, d38);
	and (d50, d15, d36);
	or (d51, d29, d31);
	nand (d52, d18, d22);
	and (d53, d7, d16);
	not (d54, d13);
	xor (d55, d12, d23);
	xor (d56, d21, d27);
	and (d57, d13, d28);
	nand (d58, d19, d34);
	and (d59, d17, d23);
	nor (d60, d6, d25);
	not (d61, d8);
	and (d62, d17, d26);
	buf (d63, d36);
	nor (d64, d8, d19);
	buf (d65, d3);
	xor (d66, d10, d19);
	buf (d67, d26);
	buf (d68, x3);
	xor (d69, d39, d46);
	and (d70, d39, d58);
	buf (d71, d65);
	or (d72, d44, d60);
	and (d73, d55, d66);
	not (d74, d16);
	buf (d75, d51);
	xnor (d76, d43, d64);
	xnor (d77, d53, d65);
	and (d78, d64);
	and (d79, d57, d61);
	or (d80, d49, d50);
	and (d81, d41, d51);
	nand (d82, d57, d63);
	not (d83, d49);
	not (d84, d46);
	nor (d85, d46, d66);
	or (d86, d47, d49);
	and (d87, d52, d54);
	and (d88, d39, d41);
	xor (d89, d50, d51);
	nand (d90, d44, d58);
	not (d91, d1);
	xor (d92, d46, d62);
	and (d93, d55, d56);
	not (d94, d54);
	not (d95, d25);
	xor (d96, d48, d54);
	nand (d97, d47, d49);
	and (d98, d43, d66);
	buf (d99, d2);
	or (d100, d56, d64);
	xor (d101, d47, d65);
	nor (d102, d43, d62);
	and (d103, d42, d60);
	xnor (d104, d46, d48);
	nor (d105, d41, d59);
	nor (d106, d42, d47);
	xor (d107, d47, d60);
	nand (d108, d59, d64);
	xor (d109, d57, d65);
	buf (d110, d6);
	nand (d111, d47, d64);
	not (d112, d50);
	not (d113, d63);
	xor (d114, d52, d54);
	not (d115, d58);
	not (d116, d64);
	or (d117, d42, d57);
	xor (d118, d66);
	and (d119, d39, d62);
	not (d120, d18);
	xnor (d121, d50, d55);
	xor (d122, d51, d54);
	xnor (d123, d46, d52);
	and (d124, d52, d58);
	xnor (d125, d39, d65);
	nor (d126, d50, d67);
	xnor (d127, d52, d58);
	nor (d128, d42, d48);
	or (d129, d46, d63);
	xnor (d130, d49);
	xor (d131, d39, d55);
	not (d132, d48);
	or (d133, d41, d66);
	or (d134, d52, d53);
	nand (d135, d62, d67);
	not (d136, d57);
	buf (d137, d57);
	buf (d138, d125);
	buf (d139, d96);
	or (d140, d96, d103);
	not (d141, d22);
	not (d142, d69);
	buf (d143, d52);
	and (d144, d138, d139);
	xor (d145, d139, d140);
	or (d146, d138, d139);
	not (d147, d97);
	and (d148, d138);
	xor (d149, d139, d140);
	nor (d150, d138, d139);
	and (d151, d139, d140);
	not (d152, d124);
	xor (d153, d139);
	buf (d154, d48);
	and (d155, d139, d140);
	or (d156, d140);
	xnor (d157, d139, d140);
	nand (d158, d139);
	or (d159, d138, d140);
	xor (d160, d140);
	xor (d161, d138, d139);
	buf (d162, d19);
	xnor (d163, d138);
	xnor (d164, d138, d140);
	xor (d165, d138, d139);
	buf (d166, d93);
	not (d167, d68);
	or (d168, d139, d140);
	buf (d169, d90);
	nand (d170, d138);
	buf (d171, d67);
	nand (d172, d139, d140);
	nor (d173, d138, d140);
	nand (d174, d138, d140);
	buf (d175, d108);
	buf (d176, d12);
	xnor (d177, d140);
	not (d178, d120);
	xor (d179, d138);
	not (d180, d36);
	nor (d181, d139);
	nor (d182, d140);
	xnor (d183, d139, d140);
	buf (d184, d137);
	nand (d185, d138, d140);
	xor (d186, d138, d140);
	and (d187, d138, d140);
	nand (d188, d139, d140);
	xnor (d189, d138, d139);
	nor (d190, d138, d139);
	nand (d191, d138, d139);
	or (d192, d138, d139);
	not (d193, d40);
	xnor (d194, d138, d140);
	not (d195, d38);
	or (d196, d138, d140);
	nand (d197, d140);
	not (d198, d129);
	not (d199, d132);
	and (d200, d154, d159);
	or (d201, d152, d175);
	nor (d202, d157, d169);
	xor (d203, d168, d194);
	xnor (d204, d155, d171);
	and (d205, d159, d162);
	xnor (d206, d169, d179);
	xor (d207, d147, d190);
	xor (d208, d150, d173);
	nand (d209, d171, d199);
	buf (d210, d104);
	not (d211, d90);
	not (d212, d146);
	and (d213, d141, d160);
	xnor (d214, d148, d188);
	nor (d215, d156, d162);
	and (d216, d162, d186);
	and (d217, d185, d187);
	nor (d218, d190, d195);
	and (d219, d189, d193);
	not (d220, d178);
	nor (d221, d161, d194);
	xor (d222, d149, d182);
	or (d223, d150, d157);
	or (d224, d147, d173);
	and (d225, d173, d190);
	not (d226, d42);
	nand (d227, d168, d191);
	nand (d228, d153, d181);
	or (d229, d157, d186);
	nand (d230, d172, d178);
	buf (d231, d102);
	buf (d232, d78);
	or (d233, d147, d194);
	and (d234, d142, d173);
	or (d235, d163, d176);
	not (d236, d95);
	buf (d237, d43);
	nor (d238, d169, d196);
	not (d239, d135);
	not (d240, d161);
	and (d241, d183, d192);
	xnor (d242, d167, d192);
	nor (d243, d150, d181);
	and (d244, d148, d188);
	and (d245, d148);
	xnor (d246, d155, d182);
	buf (d247, d198);
	or (d248, d162, d182);
	nand (d249, d141, d149);
	xnor (d250, d147, d182);
	and (d251, d145, d191);
	xor (d252, d188, d193);
	buf (d253, d21);
	nor (d254, d179, d181);
	buf (d255, d85);
	nor (d256, d176, d183);
	or (d257, d148, d166);
	or (d258, d168, d180);
	buf (d259, d167);
	nand (d260, d153, d168);
	buf (d261, d183);
	nor (d262, d150, d169);
	xor (d263, d141, d158);
	xor (d264, d147, d159);
	and (d265, d147, d156);
	xor (d266, d163, d190);
	and (d267, d144, d179);
	not (d268, d189);
	nand (d269, d155);
	and (d270, d151, d159);
	or (d271, d191);
	buf (d272, d166);
	nor (d273, d152, d187);
	buf (d274, d47);
	and (d275, d149, d177);
	or (d276, d151, d180);
	nor (d277, d144, d171);
	xnor (d278, d154, d161);
	and (d279, d174, d186);
	xnor (d280, d167, d175);
	nor (d281, d156, d163);
	buf (d282, d24);
	and (d283, d266, d276);
	xor (d284, d230, d255);
	nor (d285, d236, d239);
	nand (d286, d250, d260);
	xor (d287, d219, d243);
	nor (d288, d202, d269);
	buf (d289, d276);
	nor (d290, d207, d219);
	nand (d291, d279, d282);
	nand (d292, d226, d267);
	and (d293, d241, d249);
	and (d294, d222, d253);
	buf (d295, d49);
	buf (d296, d232);
	nor (d297, d289, d291);
	nand (d298, d283, d291);
	buf (d299, d262);
	xor (d300, d283, d294);
	buf (d301, d58);
	xnor (d302, d286, d288);
	not (d303, d91);
	not (d304, d223);
	not (d305, d287);
	or (d306, d284, d287);
	xor (d307, d283, d290);
	assign f1 = d301;
	assign f2 = d303;
endmodule
