module CCGRCG56( x0, x1, x2, x3, x4, x5, x6, x7, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13 );

	input x0, x1, x2, x3, x4, x5, x6, x7;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314, d315, d316, d317, d318, d319, d320, d321, d322, d323, d324, d325, d326, d327, d328, d329, d330, d331, d332, d333, d334, d335, d336, d337, d338, d339, d340, d341, d342, d343, d344, d345, d346, d347, d348, d349, d350, d351, d352, d353, d354, d355, d356, d357, d358, d359, d360, d361, d362, d363, d364, d365, d366, d367, d368, d369, d370, d371, d372, d373, d374, d375, d376, d377, d378, d379, d380, d381, d382, d383, d384, d385, d386, d387, d388, d389, d390, d391, d392, d393, d394, d395, d396, d397, d398, d399, d400, d401, d402, d403, d404, d405, d406, d407, d408, d409, d410, d411, d412, d413, d414, d415, d416, d417, d418, d419, d420, d421, d422, d423, d424, d425, d426, d427, d428, d429, d430, d431, d432, d433, d434, d435, d436, d437, d438, d439, d440, d441, d442, d443, d444, d445, d446, d447, d448, d449, d450, d451, d452, d453, d454, d455, d456, d457, d458, d459, d460, d461, d462, d463, d464, d465, d466, d467, d468, d469, d470, d471, d472, d473, d474, d475, d476, d477, d478, d479, d480, d481, d482, d483, d484, d485, d486, d487, d488, d489, d490, d491, d492, d493, d494, d495, d496, d497, d498, d499, d500, d501, d502, d503, d504, d505, d506, d507, d508, d509, d510, d511, d512, d513, d514, d515, d516, d517, d518, d519, d520, d521, d522, d523, d524, d525, d526, d527, d528, d529, d530, d531, d532, d533, d534, d535, d536, d537, d538, d539, d540, d541, d542, d543, d544, d545, d546, d547, d548, d549, d550, d551, d552, d553, d554, d555, d556, d557, d558, d559, d560, d561, d562, d563, d564, d565, d566, d567, d568, d569, d570, d571, d572, d573, d574, d575, d576, d577, d578, d579, d580, d581, d582, d583, d584, d585, d586, d587, d588, d589, d590, d591, d592, d593, d594, d595, d596, d597, d598, d599, d600, d601, d602, d603, d604, d605, d606, d607, d608, d609, d610, d611, d612, d613, d614, d615, d616, d617, d618, d619, d620, d621, d622, d623, d624, d625, d626, d627, d628, d629, d630, d631, d632, d633, d634, d635, d636, d637, d638, d639, d640, d641, d642, d643, d644, d645, d646, d647, d648, d649, d650, d651, d652, d653, d654, d655, d656, d657, d658, d659, d660, d661, d662, d663, d664, d665, d666, d667, d668, d669, d670, d671, d672, d673, d674, d675, d676, d677, d678, d679, d680, d681, d682, d683, d684, d685, d686, d687, d688, d689, d690, d691, d692, d693, d694, d695, d696, d697, d698, d699, d700, d701, d702, d703, d704, d705, d706, d707, d708, d709, d710, d711, d712, d713, d714, d715, d716, d717, d718, d719, d720, d721, d722, d723, d724, d725, d726, d727, d728, d729, d730, d731, d732, d733, d734, d735, d736, d737, d738, d739, d740, d741, d742, d743, d744, d745, d746, d747, d748, d749, d750, d751, d752, d753, d754, d755, d756, d757, d758, d759, d760, d761, d762, d763, d764, d765, d766, d767, d768, d769, d770, d771, d772, d773, d774, d775, d776, d777, d778, d779, d780, d781, d782, d783, d784, d785, d786, d787, d788, d789, d790, d791, d792, d793, d794, d795, d796, d797, d798, d799, d800, d801, d802, d803, d804, d805, d806, d807, d808, d809, d810, d811, d812, d813, d814, d815, d816, d817, d818, d819, d820, d821, d822, d823, d824;

	nand ( d1, x2, x4);
	buf ( d2, x5);
	nand ( d3, x6);
	nor ( d4, x0, x1);
	or ( d5, x2, x3);
	xnor ( d6, x4, x7);
	nor ( d7, x1, x4);
	and ( d8, x2);
	xor ( d9, x3, x5);
	and ( d10, x0, x2);
	nand ( d11, x6, x7);
	not ( d12, x0);
	nand ( d13, x3, x7);
	xor ( d14, x4, x7);
	nor ( d15, x1, x4);
	xnor ( d16, x3, x4);
	nor ( d17, x0, x5);
	or ( d18, x0, x3);
	not ( d19, x5);
	buf ( d20, x0);
	buf ( d21, x6);
	or ( d22, x0, x5);
	nand ( d23, x0, x6);
	nor ( d24, x0, x1);
	not ( d25, x3);
	or ( d26, x2);
	xnor ( d27, x6);
	buf ( d28, x7);
	not ( d29, x6);
	or ( d30, x2, x5);
	and ( d31, x2, x5);
	xor ( d32, x1, x6);
	nand ( d33, x3, x4);
	not ( d34, x7);
	xnor ( d35, x0, x3);
	and ( d36, x5, x7);
	or ( d37, x4, x6);
	buf ( d38, x2);
	xor ( d39, x0);
	and ( d40, d32, d38);
	not ( d41, d8);
	not ( d42, x1);
	and ( d43, d7, d37);
	buf ( d44, d19);
	buf ( d45, d3);
	not ( d46, d35);
	or ( d47, d40, d42);
	xnor ( d48, d44, d45);
	buf ( d49, d23);
	not ( d50, d25);
	xnor ( d51, d41, d45);
	buf ( d52, d43);
	and ( d53, d44, d45);
	or ( d54, d41, d45);
	buf ( d55, d18);
	nor ( d56, d41, d45);
	xnor ( d57, d41, d44);
	buf ( d58, d2);
	buf ( d59, x3);
	or ( d60, d42, d45);
	nor ( d61, d41, d45);
	or ( d62, d43, d44);
	xor ( d63, d41, d43);
	nor ( d64, d40, d44);
	buf ( d65, d28);
	and ( d66, d43, d45);
	and ( d67, d40, d42);
	xnor ( d68, d40, d41);
	buf ( d69, d6);
	not ( d70, d2);
	and ( d71, d40, d41);
	and ( d72, d44, d45);
	and ( d73, d41, d43);
	nor ( d74, d44, d45);
	nor ( d75, d40, d43);
	and ( d76, d40, d44);
	buf ( d77, d11);
	and ( d78, d43);
	xor ( d79, d43, d45);
	nor ( d80, d42, d45);
	nand ( d81, d40, d44);
	xor ( d82, d40, d44);
	or ( d83, d40, d43);
	not ( d84, d4);
	or ( d85, d40, d43);
	xnor ( d86, d42, d43);
	or ( d87, d50, d57);
	nand ( d88, d54);
	not ( d89, d15);
	xor ( d90, d54, d77);
	xnor ( d91, d48, d76);
	not ( d92, d31);
	xnor ( d93, d76, d82);
	or ( d94, d61, d72);
	xor ( d95, d57, d74);
	or ( d96, d59, d62);
	nand ( d97, d72, d73);
	not ( d98, d21);
	buf ( d99, d33);
	buf ( d100, d84);
	and ( d101, d61, d72);
	xnor ( d102, d63, d85);
	xnor ( d103, d54, d79);
	buf ( d104, d69);
	nand ( d105, d60, d71);
	nor ( d106, d67, d81);
	nor ( d107, d58, d64);
	xor ( d108, d50, d76);
	buf ( d109, d72);
	and ( d110, d50, d61);
	nand ( d111, d80);
	and ( d112, d107, d109);
	and ( d113, d94, d111);
	or ( d114, d87, d107);
	nand ( d115, d91, d102);
	and ( d116, d87, d93);
	nand ( d117, d93, d106);
	or ( d118, d103, d111);
	xor ( d119, d95, d111);
	not ( d120, d14);
	nor ( d121, d98, d111);
	or ( d122, d98, d104);
	xor ( d123, d97, d105);
	and ( d124, d89, d98);
	and ( d125, d104, d110);
	or ( d126, d95, d102);
	nand ( d127, d89, d93);
	xnor ( d128, d108, d111);
	xor ( d129, d103, d111);
	nor ( d130, d92, d103);
	xnor ( d131, d94, d108);
	buf ( d132, d82);
	xor ( d133, d93, d105);
	not ( d134, d20);
	xnor ( d135, d95, d104);
	xnor ( d136, d91, d105);
	nor ( d137, d102, d106);
	xor ( d138, d95, d110);
	xnor ( d139, d94, d110);
	nor ( d140, d113, d138);
	nor ( d141, d112, d129);
	nor ( d142, d129, d134);
	buf ( d143, d108);
	nor ( d144, d124, d136);
	not ( d145, d100);
	or ( d146, d129, d133);
	not ( d147, d139);
	buf ( d148, d10);
	nand ( d149, d112, d134);
	xnor ( d150, d124, d128);
	xnor ( d151, d118, d138);
	nor ( d152, d115, d121);
	nand ( d153, d113, d124);
	or ( d154, d120, d126);
	and ( d155, d117, d120);
	nand ( d156, d123, d135);
	nand ( d157, d114, d123);
	xor ( d158, d113);
	xor ( d159, d134, d136);
	not ( d160, d138);
	nor ( d161, d121, d139);
	buf ( d162, d44);
	not ( d163, d106);
	and ( d164, d116, d133);
	nor ( d165, d112, d117);
	and ( d166, d114, d116);
	not ( d167, d136);
	and ( d168, d135, d137);
	and ( d169, d127, d129);
	nor ( d170, d112, d113);
	nand ( d171, d124, d137);
	and ( d172, d123, d134);
	xor ( d173, d124, d131);
	xnor ( d174, d114, d125);
	and ( d175, d115, d133);
	xnor ( d176, d123, d131);
	xor ( d177, d134, d137);
	buf ( d178, d138);
	xor ( d179, d115, d121);
	nor ( d180, d127, d128);
	nor ( d181, d112, d116);
	nand ( d182, d121, d126);
	and ( d183, d112, d134);
	xnor ( d184, d113, d139);
	not ( d185, d42);
	xnor ( d186, d115, d129);
	nand ( d187, d122, d134);
	or ( d188, d147, d148);
	buf ( d189, d153);
	nand ( d190, d151, d161);
	xnor ( d191, d144, d146);
	xor ( d192, d147, d157);
	xnor ( d193, d150, d161);
	or ( d194, d166, d168);
	xnor ( d195, d145, d163);
	buf ( d196, d161);
	nand ( d197, d152, d153);
	nand ( d198, d164, d173);
	xnor ( d199, d152, d155);
	xnor ( d200, d181, d186);
	or ( d201, d157, d159);
	and ( d202, d147, d152);
	nor ( d203, d167, d168);
	nor ( d204, d151, d164);
	or ( d205, d146, d161);
	buf ( d206, d73);
	nand ( d207, d154, d166);
	nand ( d208, d190, d194);
	or ( d209, d188, d200);
	nor ( d210, d201, d204);
	nor ( d211, d188, d191);
	and ( d212, d197, d201);
	buf ( d213, d195);
	buf ( d214, d197);
	xnor ( d215, d203);
	xnor ( d216, d193, d195);
	nor ( d217, d188, d198);
	not ( d218, d45);
	and ( d219, d199, d205);
	xnor ( d220, d199, d207);
	buf ( d221, x1);
	not ( d222, d142);
	or ( d223, d210, d212);
	not ( d224, d166);
	xor ( d225, d212, d217);
	nand ( d226, d214, d216);
	nor ( d227, d214, d221);
	not ( d228, d156);
	not ( d229, d151);
	and ( d230, d209, d221);
	nand ( d231, d216, d220);
	buf ( d232, d192);
	buf ( d233, d181);
	xnor ( d234, d209, d220);
	nand ( d235, d209, d219);
	xor ( d236, d212, d216);
	not ( d237, d87);
	nand ( d238, d209, d215);
	nand ( d239, d210, d216);
	nand ( d240, d216, d217);
	or ( d241, d211, d219);
	xnor ( d242, d211, d219);
	and ( d243, d210, d216);
	and ( d244, d209, d219);
	xor ( d245, d209, d215);
	not ( d246, d110);
	and ( d247, d232, d244);
	and ( d248, d233, d246);
	or ( d249, d240, d244);
	nor ( d250, d247, d249);
	xnor ( d251, d248);
	xor ( d252, d248, d249);
	xor ( d253, d247);
	or ( d254, d249);
	nand ( d255, d247, d249);
	xnor ( d256, d247, d249);
	xor ( d257, d248, d249);
	and ( d258, d247);
	not ( d259, d214);
	nor ( d260, d247);
	not ( d261, d82);
	xor ( d262, d247, d249);
	and ( d263, d248, d249);
	nor ( d264, d248);
	nand ( d265, d247, d249);
	nor ( d266, d247, d248);
	and ( d267, d247, d248);
	or ( d268, d247, d249);
	nor ( d269, d248, d249);
	or ( d270, d247);
	nand ( d271, d249);
	buf ( d272, d235);
	and ( d273, d249);
	xnor ( d274, d247, d249);
	not ( d275, d88);
	not ( d276, d191);
	and ( d277, d248, d249);
	xnor ( d278, d248, d249);
	buf ( d279, d268);
	not ( d280, d117);
	nor ( d281, d253, d276);
	xnor ( d282, d258, d267);
	or ( d283, d251, d271);
	nand ( d284, d254, d270);
	xnor ( d285, d250, d255);
	xor ( d286, d260, d276);
	buf ( d287, d75);
	or ( d288, d250, d251);
	nand ( d289, d251, d254);
	nand ( d290, d258, d270);
	buf ( d291, d22);
	xor ( d292, d253, d273);
	not ( d293, d206);
	and ( d294, d250, d272);
	and ( d295, d251, d264);
	nor ( d296, d252, d253);
	xnor ( d297, d256, d257);
	nand ( d298, d258, d263);
	nor ( d299, d263, d269);
	and ( d300, d260, d277);
	xor ( d301, d265, d278);
	or ( d302, d263, d277);
	xnor ( d303, d263, d273);
	nor ( d304, d266, d275);
	nor ( d305, d264, d266);
	nand ( d306, d254, d257);
	xor ( d307, d269, d274);
	nor ( d308, d270, d277);
	or ( d309, d254, d267);
	and ( d310, d254, d262);
	xor ( d311, d264, d272);
	and ( d312, d265, d272);
	buf ( d313, d183);
	nor ( d314, d264, d266);
	or ( d315, d254, d260);
	or ( d316, d270, d271);
	nor ( d317, d280, d316);
	nand ( d318, d285, d311);
	xnor ( d319, d306, d316);
	xnor ( d320, d303, d304);
	or ( d321, d292, d297);
	xor ( d322, d282, d314);
	buf ( d323, d51);
	xnor ( d324, d281, d312);
	nand ( d325, d284, d295);
	nor ( d326, d281, d301);
	xor ( d327, d297, d313);
	xnor ( d328, d294, d295);
	xor ( d329, d284, d315);
	nand ( d330, d301, d304);
	nor ( d331, d301, d304);
	and ( d332, d279, d280);
	nor ( d333, d298, d308);
	xnor ( d334, d281, d294);
	not ( d335, d144);
	buf ( d336, d148);
	nand ( d337, d307, d314);
	nor ( d338, d288, d289);
	nor ( d339, d306, d307);
	xor ( d340, d292, d299);
	nor ( d341, d286, d297);
	not ( d342, d52);
	buf ( d343, d15);
	xnor ( d344, d298, d313);
	nand ( d345, d283, d297);
	xor ( d346, d290, d308);
	nand ( d347, d290, d311);
	xor ( d348, d280, d296);
	buf ( d349, d65);
	not ( d350, d165);
	or ( d351, d281, d289);
	buf ( d352, d289);
	or ( d353, d279, d304);
	and ( d354, d290, d313);
	and ( d355, d301, d316);
	xor ( d356, d282, d305);
	nor ( d357, d279, d285);
	nor ( d358, d288, d308);
	and ( d359, d291, d303);
	xor ( d360, d283, d301);
	xnor ( d361, d287, d311);
	buf ( d362, d70);
	nor ( d363, d290, d303);
	buf ( d364, d134);
	and ( d365, d327, d346);
	nor ( d366, d317, d363);
	xor ( d367, d347, d360);
	buf ( d368, d269);
	or ( d369, d331, d344);
	not ( d370, d314);
	xor ( d371, d328, d360);
	xnor ( d372, d320, d358);
	nor ( d373, d334, d360);
	xor ( d374, d352, d358);
	not ( d375, d10);
	xor ( d376, d347, d357);
	or ( d377, d328, d343);
	and ( d378, d332, d345);
	nor ( d379, d334, d337);
	nand ( d380, d319, d358);
	nor ( d381, d324, d349);
	buf ( d382, d14);
	nor ( d383, d342, d347);
	not ( d384, d311);
	nor ( d385, d324, d363);
	buf ( d386, d1);
	nor ( d387, d319, d332);
	and ( d388, d329, d344);
	xnor ( d389, d338, d341);
	and ( d390, d323, d331);
	nor ( d391, d332, d337);
	xor ( d392, d345, d357);
	buf ( d393, d129);
	nand ( d394, d356, d363);
	not ( d395, d239);
	not ( d396, d193);
	not ( d397, d334);
	nor ( d398, d318, d360);
	xor ( d399, d318, d338);
	xor ( d400, d321, d348);
	buf ( d401, d184);
	not ( d402, d332);
	buf ( d403, d359);
	nor ( d404, d343, d349);
	or ( d405, d387, d394);
	xor ( d406, d372, d394);
	nand ( d407, d367, d388);
	nor ( d408, d370);
	not ( d409, d86);
	nor ( d410, d369, d379);
	and ( d411, d379, d392);
	xor ( d412, d369, d396);
	xor ( d413, d364, d376);
	xor ( d414, d375, d384);
	buf ( d415, d126);
	and ( d416, d367, d372);
	buf ( d417, d272);
	or ( d418, d375, d384);
	xor ( d419, d369, d373);
	xor ( d420, d373);
	buf ( d421, d141);
	and ( d422, d389, d397);
	or ( d423, d377, d400);
	buf ( d424, d299);
	nor ( d425, d409);
	and ( d426, d413);
	xnor ( d427, d418, d421);
	buf ( d428, d222);
	nor ( d429, d407, d408);
	buf ( d430, d39);
	nor ( d431, d405, d423);
	xor ( d432, d415, d421);
	nor ( d433, d406, d419);
	or ( d434, d411, d415);
	xor ( d435, d408, d423);
	nor ( d436, d406, d417);
	buf ( d437, d127);
	or ( d438, d414, d420);
	buf ( d439, d253);
	nand ( d440, d412, d419);
	xor ( d441, d412, d416);
	and ( d442, d412, d419);
	buf ( d443, d123);
	xor ( d444, d409, d410);
	not ( d445, d162);
	and ( d446, d408, d409);
	nor ( d447, d426, d437);
	nor ( d448, d428, d432);
	buf ( d449, d86);
	and ( d450, d428, d442);
	xnor ( d451, d438, d442);
	or ( d452, d439, d441);
	buf ( d453, d241);
	xnor ( d454, d427, d441);
	not ( d455, d324);
	or ( d456, d427, d432);
	xor ( d457, d429, d434);
	not ( d458, d432);
	xor ( d459, d453);
	and ( d460, d449, d451);
	nor ( d461, d452, d457);
	and ( d462, d452, d456);
	buf ( d463, d213);
	nand ( d464, d454, d456);
	nor ( d465, d450, d454);
	buf ( d466, d401);
	nor ( d467, d449, d455);
	not ( d468, d396);
	xor ( d469, d456);
	xnor ( d470, d447, d454);
	and ( d471, d447, d454);
	nand ( d472, d454, d457);
	nand ( d473, d453, d456);
	or ( d474, d447, d453);
	and ( d475, d448);
	xnor ( d476, d447, d449);
	nand ( d477, d455, d456);
	nor ( d478, d449, d457);
	or ( d479, d449, d450);
	xor ( d480, d453, d454);
	nor ( d481, d451, d452);
	buf ( d482, d206);
	nor ( d483, d447, d456);
	not ( d484, d129);
	xnor ( d485, d449, d450);
	xnor ( d486, d447);
	buf ( d487, d227);
	xnor ( d488, d453, d455);
	buf ( d489, d386);
	xor ( d490, d452, d453);
	not ( d491, d74);
	xor ( d492, d447, d455);
	or ( d493, d448, d452);
	not ( d494, d22);
	nor ( d495, d449, d451);
	and ( d496, d450, d455);
	nand ( d497, d447, d450);
	or ( d498, d448, d453);
	or ( d499, d447, d448);
	xnor ( d500, d450, d454);
	xor ( d501, d448, d455);
	and ( d502, d448, d455);
	buf ( d503, d4);
	xnor ( d504, d462, d483);
	and ( d505, d484, d499);
	xor ( d506, d465, d473);
	buf ( d507, d406);
	nand ( d508, d471, d480);
	and ( d509, d464, d476);
	or ( d510, d474, d493);
	nand ( d511, d462, d485);
	and ( d512, d468, d482);
	xnor ( d513, d473, d496);
	nand ( d514, d487, d497);
	xor ( d515, d463, d497);
	and ( d516, d463, d487);
	xor ( d517, d499, d501);
	not ( d518, d382);
	or ( d519, d472, d489);
	nand ( d520, d466, d467);
	xor ( d521, d458, d484);
	xnor ( d522, d464, d470);
	nor ( d523, d469, d474);
	nor ( d524, d458, d462);
	nand ( d525, d470, d486);
	xor ( d526, d477, d490);
	and ( d527, d459, d502);
	buf ( d528, d457);
	buf ( d529, d294);
	and ( d530, d458, d471);
	or ( d531, d463, d476);
	or ( d532, d469, d480);
	nand ( d533, d476, d494);
	or ( d534, d461, d494);
	or ( d535, d473, d479);
	xnor ( d536, d482, d490);
	buf ( d537, d473);
	or ( d538, d467, d484);
	not ( d539, d60);
	buf ( d540, d336);
	or ( d541, d480, d495);
	not ( d542, d449);
	nor ( d543, d462, d476);
	nand ( d544, d468, d489);
	nor ( d545, d460, d482);
	and ( d546, d464, d500);
	nor ( d547, d468, d472);
	nor ( d548, d463, d477);
	nand ( d549, d537, d548);
	nand ( d550, d545);
	not ( d551, d374);
	xnor ( d552, d535);
	nor ( d553, d522, d536);
	and ( d554, d511, d512);
	buf ( d555, d546);
	not ( d556, d9);
	not ( d557, d329);
	nand ( d558, d514, d517);
	or ( d559, d507, d527);
	nand ( d560, d510, d541);
	xnor ( d561, d531, d536);
	and ( d562, d509, d544);
	xnor ( d563, d558, d560);
	or ( d564, d554, d555);
	xnor ( d565, d550, d557);
	not ( d566, d428);
	or ( d567, d555);
	nand ( d568, d549, d559);
	xor ( d569, d565, d566);
	nand ( d570, d563);
	xor ( d571, d567, d568);
	xor ( d572, d566, d568);
	and ( d573, d564, d568);
	or ( d574, d566, d568);
	and ( d575, d565, d566);
	or ( d576, d564, d566);
	nand ( d577, d565, d566);
	buf ( d578, d246);
	buf ( d579, d393);
	xor ( d580, d564, d566);
	nor ( d581, d566, d567);
	not ( d582, d326);
	nor ( d583, d563, d564);
	nor ( d584, d566);
	nand ( d585, d564, d566);
	buf ( d586, d92);
	buf ( d587, d377);
	nand ( d588, d567, d568);
	not ( d589, d439);
	buf ( d590, d562);
	and ( d591, d576, d589);
	not ( d592, d221);
	buf ( d593, d322);
	nand ( d594, d572, d575);
	and ( d595, d573, d589);
	xor ( d596, d575, d580);
	or ( d597, d571, d590);
	xnor ( d598, d570);
	nor ( d599, d587, d589);
	xnor ( d600, d570, d578);
	or ( d601, d587, d590);
	buf ( d602, d531);
	or ( d603, d573, d589);
	xnor ( d604, d577, d588);
	not ( d605, d51);
	or ( d606, d579, d587);
	xnor ( d607, d577, d583);
	buf ( d608, d525);
	or ( d609, d578);
	and ( d610, d578, d590);
	buf ( d611, d349);
	not ( d612, d534);
	xnor ( d613, d578, d587);
	xnor ( d614, d575, d588);
	xnor ( d615, d571, d585);
	nand ( d616, d572, d581);
	nand ( d617, d571, d578);
	xor ( d618, d583, d586);
	or ( d619, d582, d585);
	xnor ( d620, d582, d590);
	buf ( d621, d58);
	nand ( d622, d580, d581);
	buf ( d623, d311);
	and ( d624, d570, d571);
	and ( d625, d571, d581);
	or ( d626, d582, d583);
	nand ( d627, d581, d584);
	xor ( d628, d569, d570);
	xnor ( d629, d574, d587);
	or ( d630, d586, d588);
	nor ( d631, d576, d578);
	nand ( d632, d574, d588);
	or ( d633, d574, d583);
	nor ( d634, d578, d579);
	xnor ( d635, d580, d588);
	not ( d636, d33);
	xor ( d637, d596, d603);
	xnor ( d638, d613, d622);
	nand ( d639, d604, d618);
	xor ( d640, d597, d619);
	buf ( d641, d102);
	or ( d642, d593, d616);
	nand ( d643, d620, d624);
	and ( d644, d594, d602);
	buf ( d645, d199);
	or ( d646, d593, d614);
	or ( d647, d608, d634);
	and ( d648, d608, d620);
	and ( d649, d611, d612);
	xnor ( d650, d608, d630);
	nand ( d651, d626, d633);
	xor ( d652, d604, d619);
	buf ( d653, d506);
	nand ( d654, d612, d634);
	nand ( d655, d601, d630);
	or ( d656, d601, d607);
	not ( d657, d225);
	xnor ( d658, d599, d602);
	nand ( d659, d613, d618);
	nand ( d660, d609, d614);
	xor ( d661, d649, d652);
	nor ( d662, d636, d644);
	buf ( d663, d445);
	or ( d664, d643, d651);
	not ( d665, d361);
	xor ( d666, d638, d641);
	nand ( d667, d650, d658);
	or ( d668, d648, d658);
	nand ( d669, d636, d650);
	nor ( d670, d642, d659);
	buf ( d671, d53);
	nor ( d672, d646, d649);
	nor ( d673, d644, d654);
	or ( d674, d637, d646);
	and ( d675, d639, d644);
	nand ( d676, d638, d652);
	nand ( d677, d642, d654);
	xnor ( d678, d640, d643);
	nor ( d679, d646, d654);
	nor ( d680, d653, d656);
	xor ( d681, d638, d654);
	xnor ( d682, d648, d655);
	nor ( d683, d645, d650);
	or ( d684, d637, d638);
	and ( d685, d637, d650);
	xnor ( d686, d636, d649);
	xnor ( d687, d636, d658);
	xor ( d688, d649, d651);
	buf ( d689, d403);
	xnor ( d690, d649, d660);
	and ( d691, d650, d657);
	and ( d692, d650, d659);
	buf ( d693, d7);
	or ( d694, d653, d655);
	nor ( d695, d643, d658);
	xnor ( d696, d655, d660);
	nand ( d697, d649);
	and ( d698, d642, d645);
	not ( d699, d560);
	nand ( d700, d642, d654);
	nor ( d701, d653, d660);
	nand ( d702, d666, d677);
	nor ( d703, d662, d666);
	nand ( d704, d694, d696);
	nand ( d705, d668, d680);
	nand ( d706, d677, d681);
	nand ( d707, d688, d700);
	xor ( d708, d682, d686);
	nor ( d709, d669, d698);
	buf ( d710, d700);
	not ( d711, d167);
	nand ( d712, d668, d681);
	nor ( d713, d667, d674);
	nand ( d714, d677, d687);
	and ( d715, d663, d677);
	nand ( d716, d680, d682);
	not ( d717, d186);
	or ( d718, d682, d683);
	not ( d719, d201);
	buf ( d720, d532);
	nor ( d721, d662, d678);
	xor ( d722, d677);
	xnor ( d723, d690, d694);
	nor ( d724, d671, d673);
	xor ( d725, d669, d697);
	buf ( d726, d88);
	or ( d727, d679, d680);
	or ( d728, d680, d690);
	xnor ( d729, d676, d694);
	or ( d730, d690, d701);
	not ( d731, d688);
	nand ( d732, d661, d669);
	xnor ( d733, d674, d676);
	or ( d734, d671, d676);
	and ( d735, d665, d668);
	xnor ( d736, d675, d688);
	xnor ( d737, d682, d694);
	nor ( d738, d673, d678);
	not ( d739, d37);
	and ( d740, d686, d687);
	or ( d741, d662, d669);
	buf ( d742, d411);
	buf ( d743, d519);
	or ( d744, d711, d724);
	xnor ( d745, d716, d719);
	nand ( d746, d711, d723);
	xor ( d747, d703, d737);
	or ( d748, d717, d733);
	not ( d749, d429);
	xnor ( d750, d721, d743);
	nor ( d751, d711, d736);
	xor ( d752, d720, d735);
	xnor ( d753, d717, d730);
	nand ( d754, d722, d739);
	not ( d755, d150);
	xor ( d756, d724, d741);
	not ( d757, d554);
	buf ( d758, d621);
	xor ( d759, d708, d719);
	buf ( d760, d217);
	not ( d761, d441);
	not ( d762, d253);
	buf ( d763, d480);
	and ( d764, d702, d704);
	not ( d765, d666);
	nor ( d766, d705, d720);
	and ( d767, d704, d724);
	buf ( d768, d559);
	or ( d769, d713, d730);
	xnor ( d770, d716, d728);
	or ( d771, d722, d723);
	nor ( d772, d706, d720);
	nand ( d773, d713, d730);
	and ( d774, d702, d719);
	and ( d775, d758, d761);
	not ( d776, d352);
	not ( d777, d304);
	xor ( d778, d758, d774);
	nor ( d779, d750, d770);
	and ( d780, d747, d764);
	buf ( d781, d52);
	not ( d782, d49);
	not ( d783, d77);
	not ( d784, d46);
	nand ( d785, d759, d769);
	xnor ( d786, d762, d771);
	nand ( d787, d760, d761);
	xnor ( d788, d778, d782);
	nand ( d789, d777, d782);
	and ( d790, d777, d780);
	xnor ( d791, d785);
	xor ( d792, d786);
	or ( d793, d775, d781);
	xor ( d794, d777, d786);
	xnor ( d795, d781, d785);
	nand ( d796, d778);
	and ( d797, d786, d787);
	or ( d798, d779);
	and ( d799, d780, d785);
	nor ( d800, d780, d781);
	nor ( d801, d783, d785);
	buf ( d802, d224);
	xor ( d803, d780, d784);
	xnor ( d804, d778, d780);
	nand ( d805, d781, d787);
	or ( d806, d779, d787);
	or ( d807, d781, d787);
	buf ( d808, d783);
	xnor ( d809, d785, d786);
	not ( d810, d381);
	or ( d811, d782, d787);
	and ( d812, d783, d787);
	or ( d813, d777, d781);
	or ( d814, d777, d787);
	nor ( d815, d777, d780);
	nand ( d816, d776, d782);
	buf ( d817, d431);
	not ( d818, d384);
	or ( d819, d782, d783);
	or ( d820, d779, d784);
	or ( d821, d777, d781);
	buf ( d822, d307);
	xnor ( d823, d779, d782);
	xor ( d824, d776, d777);
	assign f1 = d811;
	assign f2 = d814;
	assign f3 = d807;
	assign f4 = d809;
	assign f5 = d823;
	assign f6 = d807;
	assign f7 = d824;
	assign f8 = d798;
	assign f9 = d818;
	assign f10 = d801;
	assign f11 = d792;
	assign f12 = d811;
	assign f13 = d798;
endmodule
