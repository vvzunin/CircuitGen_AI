module CCGRCG59( x0, x1, x2, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12 );

	input x0, x1, x2;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121;

	or (d1, x0);
	buf (d2, x2);
	nor (d3, x0, x1);
	nor (d4, x0, x2);
	nor (d5, x2);
	buf (d6, x0);
	xnor (d7, x0, x2);
	nor (d8, x0, x1);
	or (d9, x1, x2);
	and (d10, x0);
	and (d11, x0, x2);
	or (d12, d4, d11);
	nand (d13, d8, d9);
	nor (d14, d3, d6);
	not (d15, d9);
	xor (d16, d7, d10);
	xnor (d17, d5, d6);
	and (d18, d5, d11);
	nor (d19, d7, d11);
	nor (d20, d6, d10);
	xor (d21, d1, d5);
	xor (d22, d1, d10);
	and (d23, d1, d3);
	xor (d24, d1, d8);
	nor (d25, d3, d4);
	nand (d26, d2, d6);
	xor (d27, d2, d7);
	nor (d28, d10);
	nand (d29, d8, d10);
	xor (d30, d3, d10);
	not (d31, d5);
	buf (d32, d11);
	not (d33, d1);
	not (d34, x2);
	not (d35, d27);
	xor (d36, d22, d23);
	nor (d37, d22, d26);
	xor (d38, d23, d32);
	and (d39, d25, d31);
	xnor (d40, d30, d33);
	xor (d41, d14, d30);
	buf (d42, d2);
	buf (d43, d26);
	not (d44, d26);
	xor (d45, d20, d34);
	xnor (d46, d34);
	nor (d47, d31, d33);
	nor (d48, d13, d15);
	buf (d49, d3);
	or (d50, d22, d26);
	or (d51, d12, d27);
	not (d52, d21);
	xnor (d53, d13, d27);
	or (d54, d15, d17);
	or (d55, d17, d30);
	xor (d56, d18, d24);
	not (d57, d7);
	xor (d58, d12, d14);
	xor (d59, d27);
	xor (d60, d40, d57);
	buf (d61, d41);
	buf (d62, d40);
	not (d63, d52);
	nor (d64, d50, d56);
	not (d65, d28);
	not (d66, d44);
	nor (d67, d46, d52);
	or (d68, d41, d46);
	xnor (d69, d44, d51);
	xnor (d70, d39, d54);
	buf (d71, d47);
	xnor (d72, d36, d54);
	or (d73, d41, d51);
	nor (d74, d39, d54);
	nand (d75, d45, d47);
	nor (d76, d39, d46);
	nor (d77, d70, d72);
	xor (d78, d76);
	nor (d79, d70, d75);
	not (d80, d13);
	xnor (d81, d67, d73);
	or (d82, d73);
	and (d83, d61, d73);
	xor (d84, d71, d73);
	not (d85, d12);
	nand (d86, d65, d72);
	nand (d87, d66, d73);
	and (d88, d65, d66);
	nor (d89, d65, d76);
	nand (d90, d72, d76);
	nand (d91, d70, d72);
	not (d92, d60);
	nor (d93, d70, d75);
	or (d94, d65, d69);
	xor (d95, d64, d67);
	xnor (d96, d60, d66);
	nor (d97, d67, d69);
	buf (d98, d13);
	or (d99, d60, d65);
	xor (d100, d69);
	nor (d101, d62, d66);
	or (d102, d61, d72);
	nor (d103, d64, d70);
	xnor (d104, d64, d70);
	nand (d105, d64, d65);
	not (d106, d51);
	buf (d107, d60);
	xnor (d108, d61, d66);
	or (d109, d65);
	nand (d110, d62, d68);
	or (d111, d68, d69);
	or (d112, d67, d71);
	xor (d113, d66, d70);
	buf (d114, d29);
	not (d115, d40);
	xor (d116, d66, d67);
	and (d117, d62, d73);
	nor (d118, d73, d74);
	and (d119, d64, d69);
	nand (d120, d69, d72);
	buf (d121, d23);
	assign f1 = d121;
	assign f2 = d88;
	assign f3 = d101;
	assign f4 = d83;
	assign f5 = d93;
	assign f6 = d120;
	assign f7 = d119;
	assign f8 = d87;
	assign f9 = d85;
	assign f10 = d118;
	assign f11 = d105;
	assign f12 = d104;
endmodule
