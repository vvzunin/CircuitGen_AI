module CCGRCG8( x0, x1, f1, f2, f3, f4, f5, f6 );

	input x0, x1;
	output f1, f2, f3, f4, f5, f6;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106;

	not (d1, x0);
	and (d2, x0, x1);
	xor (d3, x0);
	or (d4, x0, x1);
	and (d5, x0, x1);
	nor (d6, x1);
	buf (d7, x0);
	not (d8, x1);
	xor (d9, x0, x1);
	xor (d10, x1);
	xnor (d11, x0, x1);
	nor (d12, x0, x1);
	nand (d13, x1);
	xnor (d14, x0, x1);
	nor (d15, x0, x1);
	or (d16, x0);
	xor (d17, x0, x1);
	xor (d18, d8, d9);
	and (d19, d2, d7);
	xor (d20, d10, d12);
	xor (d21, d11, d14);
	buf (d22, d3);
	not (d23, d5);
	xnor (d24, d12, d14);
	nor (d25, d10, d13);
	not (d26, d7);
	xor (d27, d1, d3);
	nor (d28, d10, d14);
	xor (d29, d2, d15);
	xnor (d30, d10, d15);
	not (d31, d13);
	and (d32, d4, d17);
	nand (d33, d6, d10);
	or (d34, d8, d9);
	and (d35, d2, d9);
	and (d36, d10, d17);
	or (d37, d10, d12);
	nor (d38, d13, d16);
	and (d39, d2, d13);
	xnor (d40, d5, d8);
	xnor (d41, d2, d4);
	xor (d42, d3, d9);
	xor (d43, d5, d13);
	and (d44, d8, d13);
	not (d45, d11);
	nand (d46, d12, d17);
	or (d47, d11, d14);
	not (d48, d14);
	and (d49, d1, d7);
	xor (d50, d4, d14);
	or (d51, d12, d15);
	xor (d52, d1, d14);
	buf (d53, d1);
	nand (d54, d49, d50);
	nor (d55, d44, d47);
	nand (d56, d25, d29);
	nor (d57, d44, d51);
	nor (d58, d40, d50);
	xor (d59, d29, d37);
	xor (d60, d28, d37);
	xnor (d61, d41, d49);
	xor (d62, d47, d49);
	or (d63, d24, d41);
	not (d64, d15);
	buf (d65, d19);
	not (d66, d52);
	and (d67, d20, d30);
	or (d68, d42, d44);
	xnor (d69, d24, d32);
	xnor (d70, d29);
	buf (d71, d31);
	nand (d72, d55, d60);
	buf (d73, d33);
	buf (d74, d17);
	xnor (d75, d56, d60);
	and (d76, d54, d68);
	xnor (d77, d55, d62);
	xnor (d78, d54, d58);
	not (d79, d51);
	and (d80, d67, d70);
	or (d81, d57, d59);
	or (d82, d56, d71);
	and (d83, d62, d66);
	xnor (d84, d64, d71);
	xor (d85, d57, d60);
	xnor (d86, d55, d70);
	xor (d87, d56, d69);
	and (d88, d62, d69);
	or (d89, d65, d68);
	buf (d90, d63);
	xor (d91, d70, d71);
	nor (d92, d59, d71);
	nand (d93, d61, d69);
	or (d94, d62, d70);
	and (d95, d68);
	not (d96, d42);
	nand (d97, d54, d60);
	nand (d98, d61, d63);
	and (d99, d66, d68);
	nand (d100, d64, d70);
	nor (d101, d57, d71);
	buf (d102, d49);
	not (d103, d21);
	buf (d104, d28);
	or (d105, d60, d67);
	or (d106, d55, d56);
	assign f1 = d83;
	assign f2 = d86;
	assign f3 = d92;
	assign f4 = d106;
	assign f5 = d77;
	assign f6 = d93;
endmodule
