module CCGRCG186( x0, x1, x2, x3, x4, x5, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17, f18, f19 );

	input x0, x1, x2, x3, x4, x5;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17, f18, f19;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63;

	buf (d1, x3);
	xor (d2, x2, x3);
	nor (d3, x0, x3);
	or (d4, x0, x4);
	nand (d5, x0);
	nor (d6, x0, x4);
	xor (d7, x3, x5);
	xnor (d8, x0, x2);
	xnor (d9, x0, x4);
	nor (d10, x1);
	xnor (d11, x3, x5);
	or (d12, x3);
	nand (d13, x1, x4);
	xor (d14, x0, x4);
	or (d15, x1, x4);
	buf (d16, x0);
	buf (d17, x1);
	and (d18, x1, x4);
	and (d19, x3, x5);
	and (d20, x4, x5);
	buf (d21, x5);
	or (d22, x1, x3);
	buf (d23, x2);
	not (d24, x5);
	xnor (d25, x2, x5);
	xor (d26, x0, x3);
	nand (d27, x0, x2);
	buf (d28, x4);
	xor (d29, x1, x2);
	xnor (d30, x2, x5);
	nand (d31, x2, x5);
	nand (d32, x0, x4);
	xnor (d33, x0, x2);
	xnor (d34, x1, x5);
	and (d35, x0);
	and (d36, x1, x4);
	or (d37, x3, x4);
	xor (d38, x3);
	nor (d39, x0, x1);
	xor (d40, x3, x5);
	and (d41, x3);
	nor (d42, x2, x5);
	nand (d43, x4, x5);
	nand (d44, x0, x5);
	not (d45, x4);
	nand (d46, x0, x1);
	nand (d47, x1, x5);
	xor (d48, x1);
	nor (d49, x2);
	or (d50, x5);
	xor (d51, x2, x5);
	nand (d52, x3, x5);
	not (d53, x0);
	not (d54, d38);
	nor (d55, d21, d33);
	and (d56, d21, d50);
	xor (d57, d2, d15);
	or (d58, d44, d48);
	xor (d59, d3, d44);
	nor (d60, d18, d48);
	and (d61, d40, d46);
	or (d62, d33, d50);
	xor (d63, d15, d34);
	assign f1 = d62;
	assign f2 = d54;
	assign f3 = d59;
	assign f4 = d60;
	assign f5 = d60;
	assign f6 = d63;
	assign f7 = d55;
	assign f8 = d63;
	assign f9 = d63;
	assign f10 = d57;
	assign f11 = d62;
	assign f12 = d58;
	assign f13 = d57;
	assign f14 = d61;
	assign f15 = d59;
	assign f16 = d62;
	assign f17 = d63;
	assign f18 = d55;
	assign f19 = d55;
endmodule
