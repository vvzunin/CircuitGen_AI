module CCGRCG38( x0, x1, x2, f1, f2 );

	input x0, x1, x2;
	output f1, f2;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142;

	xor (d1, x1, x2);
	or (d2, x0, x2);
	not (d3, x0);
	xnor (d4, x0, x2);
	nand (d5, x1, x2);
	and (d6, x1, x2);
	buf (d7, x1);
	not (d8, x1);
	xor (d9, x0, x1);
	xor (d10, x2);
	or (d11, x1, x2);
	xnor (d12, x1);
	and (d13, x0, x1);
	nor (d14, x0, x2);
	xor (d15, x0, x2);
	or (d16, x1);
	xnor (d17, x2);
	nor (d18, x0);
	nor (d19, x1);
	xnor (d20, x0);
	xnor (d21, x0, x2);
	and (d22, x0, x1);
	xor (d23, x1);
	buf (d24, x0);
	and (d25, x1);
	nand (d26, x0, x2);
	nand (d27, x0, x1);
	nand (d28, x1);
	nor (d29, x0, x2);
	and (d30, x1, x2);
	and (d31, x0, x2);
	xnor (d32, x0, x1);
	or (d33, x1, x2);
	nand (d34, x2);
	buf (d35, x2);
	not (d36, x2);
	or (d37, x2);
	nor (d38, x1, x2);
	nand (d39, x0);
	nor (d40, x0, x1);
	nor (d41, x0, x1);
	nor (d42, x2);
	xnor (d43, x1, x2);
	or (d44, x0, x1);
	xor (d45, x1, x2);
	or (d46, x0, x1);
	xnor (d47, x0, x1);
	or (d48, x0);
	nand (d49, x0, x2);
	and (d50, x0, x2);
	buf (d51, d1);
	nand (d52, d10, d21);
	xnor (d53, d7, d48);
	xnor (d54, d8);
	xnor (d55, d12, d26);
	buf (d56, d7);
	buf (d57, d6);
	nand (d58, d13, d14);
	nand (d59, d41, d49);
	not (d60, d6);
	nor (d61, d12, d46);
	and (d62, d9, d17);
	nand (d63, d29, d32);
	buf (d64, d26);
	or (d65, d19, d46);
	and (d66, d32, d41);
	xnor (d67, d25, d33);
	xor (d68, d3, d18);
	or (d69, d13);
	not (d70, d24);
	not (d71, d36);
	xor (d72, d31, d32);
	xnor (d73, d6, d19);
	and (d74, d3, d44);
	xnor (d75, d31, d36);
	and (d76, d23);
	nand (d77, d3, d15);
	nand (d78, d22, d47);
	xor (d79, d22, d23);
	or (d80, d18, d39);
	or (d81, d14, d23);
	xor (d82, d19, d28);
	nor (d83, d13, d35);
	not (d84, d14);
	not (d85, d20);
	xnor (d86, d25, d27);
	xnor (d87, d33, d49);
	not (d88, d37);
	xnor (d89, d7, d40);
	xnor (d90, d5, d42);
	or (d91, d15, d25);
	xnor (d92, d10, d42);
	or (d93, d3, d43);
	xor (d94, d9, d35);
	xor (d95, d21, d25);
	not (d96, d47);
	and (d97, d10, d39);
	and (d98, d12, d36);
	nor (d99, d13, d31);
	not (d100, d5);
	and (d101, d44, d48);
	xor (d102, d28, d42);
	and (d103, d6, d26);
	xor (d104, d1, d48);
	and (d105, d14, d29);
	xnor (d106, d3, d46);
	xnor (d107, d44, d50);
	nor (d108, d6, d12);
	or (d109, d3, d41);
	xnor (d110, d17, d32);
	buf (d111, d27);
	not (d112, d1);
	xor (d113, d22, d40);
	and (d114, d4, d47);
	xor (d115, d23, d28);
	nor (d116, d14, d41);
	nand (d117, d11, d48);
	or (d118, d18, d36);
	xnor (d119, d36, d48);
	nand (d120, d8, d21);
	and (d121, d17, d21);
	not (d122, d25);
	xor (d123, d5, d28);
	xnor (d124, d10, d41);
	xor (d125, d3, d49);
	or (d126, d18, d41);
	nand (d127, d14, d29);
	or (d128, d17, d45);
	and (d129, d6, d38);
	nand (d130, d12, d21);
	xnor (d131, d9, d42);
	and (d132, d13, d25);
	xnor (d133, d19, d21);
	xnor (d134, d5, d38);
	buf (d135, d38);
	nor (d136, d7, d24);
	xnor (d137, d35, d38);
	nand (d138, d7, d48);
	not (d139, d27);
	xor (d140, d28, d47);
	buf (d141, d11);
	xor (d142, d27, d40);
	assign f1 = d62;
	assign f2 = d98;
endmodule
