module CCGRCG173( x0, x1, x2, x3, x4, x5, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12 );

	input x0, x1, x2, x3, x4, x5;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314, d315, d316, d317, d318, d319, d320, d321, d322, d323, d324, d325, d326, d327, d328, d329, d330, d331, d332, d333, d334, d335, d336, d337, d338, d339, d340, d341, d342, d343, d344, d345, d346, d347, d348, d349, d350, d351, d352, d353, d354, d355, d356, d357, d358, d359, d360, d361, d362, d363, d364, d365, d366, d367, d368, d369, d370, d371, d372, d373, d374, d375, d376, d377, d378, d379, d380, d381, d382, d383, d384, d385, d386, d387, d388, d389, d390, d391, d392, d393, d394, d395, d396, d397, d398, d399, d400, d401, d402, d403, d404, d405, d406, d407, d408, d409, d410, d411, d412, d413, d414, d415, d416, d417, d418, d419, d420, d421, d422, d423, d424, d425, d426, d427, d428, d429, d430, d431, d432, d433, d434, d435, d436, d437, d438, d439, d440, d441, d442, d443, d444, d445, d446, d447, d448, d449, d450, d451, d452, d453, d454, d455, d456, d457, d458, d459, d460, d461, d462, d463, d464, d465, d466, d467, d468, d469, d470, d471, d472, d473, d474, d475, d476, d477, d478, d479, d480, d481, d482, d483, d484, d485, d486, d487, d488, d489, d490, d491, d492, d493, d494, d495, d496, d497, d498, d499, d500, d501, d502, d503, d504, d505, d506, d507, d508, d509, d510, d511, d512, d513, d514, d515, d516, d517, d518, d519, d520, d521, d522, d523, d524, d525, d526, d527, d528, d529, d530, d531, d532, d533, d534, d535, d536, d537, d538, d539, d540, d541, d542, d543, d544, d545, d546, d547, d548, d549, d550, d551, d552, d553, d554, d555, d556, d557, d558, d559, d560, d561, d562, d563, d564, d565, d566, d567, d568, d569, d570, d571, d572, d573, d574, d575, d576, d577, d578, d579, d580, d581, d582, d583, d584, d585;

	xnor (d1, x0, x3);
	and (d2, x1, x2);
	nor (d3, x1);
	xnor (d4, x0, x2);
	xnor (d5, x4, x5);
	and (d6, x2, x5);
	not (d7, x2);
	xor (d8, x3);
	xor (d9, x4, x5);
	xor (d10, x2);
	or (d11, x1, x2);
	nand (d12, x2, x3);
	and (d13, x3, x5);
	xor (d14, x1, x2);
	nand (d15, x0, x2);
	xor (d16, x1, x3);
	nor (d17, x2, x3);
	xor (d18, x1, x2);
	and (d19, x2, x3);
	or (d20, x3);
	nand (d21, x3, x5);
	not (d22, x0);
	nand (d23, x1, x2);
	nand (d24, x0, x3);
	buf (d25, x3);
	xnor (d26, x1);
	xor (d27, x1, x4);
	not (d28, x4);
	nand (d29, x2, x4);
	and (d30, x2, x5);
	or (d31, x1, x4);
	not (d32, x3);
	or (d33, x2, x5);
	and (d34, x1, x2);
	or (d35, x0, x4);
	or (d36, x5);
	xnor (d37, x1, x4);
	or (d38, x1, x3);
	or (d39, x1, x5);
	nor (d40, x0, x3);
	nand (d41, x0);
	nor (d42, x4);
	xnor (d43, x3, x5);
	buf (d44, x2);
	and (d45, x1, x3);
	not (d46, x5);
	and (d47, x3, x5);
	and (d48, x0, x1);
	xor (d49, x2, x3);
	and (d50, x0);
	buf (d51, x4);
	or (d52, x2, x5);
	or (d53, x0, x2);
	xor (d54, x2, x5);
	buf (d55, x1);
	xnor (d56, x3);
	and (d57, x1);
	nor (d58, x0, x5);
	nand (d59, x2, x5);
	xor (d60, x1, x5);
	nand (d61, x3, x4);
	buf (d62, x0);
	xnor (d63, x0, x2);
	and (d64, x0, x3);
	xnor (d65, d13, d16);
	or (d66, d40, d47);
	or (d67, d4, d39);
	nand (d68, d20, d53);
	or (d69, d31, d32);
	nor (d70, d46, d47);
	and (d71, d11, d42);
	nand (d72, d3, d9);
	xor (d73, d1, d41);
	or (d74, d11, d34);
	buf (d75, d57);
	and (d76, d6, d56);
	nor (d77, d18, d33);
	not (d78, d54);
	buf (d79, d58);
	nand (d80, d10, d35);
	or (d81, d34, d46);
	not (d82, d3);
	not (d83, d29);
	nand (d84, d3, d36);
	nor (d85, d21, d49);
	nand (d86, d50, d54);
	not (d87, d52);
	xor (d88, d58, d61);
	buf (d89, d7);
	nand (d90, d2, d50);
	xnor (d91, d47, d63);
	xnor (d92, d4, d57);
	nand (d93, d5, d62);
	xor (d94, d5, d44);
	xnor (d95, d16, d36);
	nand (d96, d4, d34);
	and (d97, d19, d64);
	nand (d98, d39, d57);
	or (d99, d39, d42);
	or (d100, d29, d31);
	buf (d101, d47);
	and (d102, d7, d19);
	nor (d103, d38, d41);
	buf (d104, d14);
	xnor (d105, d3, d23);
	nor (d106, d23, d41);
	not (d107, d49);
	xor (d108, d9, d10);
	and (d109, d15, d22);
	nand (d110, d41, d47);
	not (d111, d43);
	xnor (d112, d1, d13);
	nand (d113, d12, d56);
	not (d114, d44);
	buf (d115, d22);
	and (d116, d5, d22);
	xnor (d117, d44);
	nand (d118, d2, d47);
	buf (d119, d32);
	not (d120, d16);
	nor (d121, d26, d34);
	not (d122, d19);
	nand (d123, d21, d37);
	xnor (d124, d46, d59);
	nand (d125, d17, d33);
	and (d126, d50);
	not (d127, d28);
	and (d128, d28, d47);
	not (d129, d62);
	xor (d130, d24, d55);
	not (d131, d56);
	xor (d132, d35, d40);
	and (d133, d28, d29);
	xor (d134, d15, d27);
	buf (d135, d42);
	nor (d136, d22, d38);
	buf (d137, d60);
	xnor (d138, d73, d111);
	xor (d139, d100, d105);
	or (d140, d74, d101);
	xnor (d141, d136, d137);
	and (d142, d77, d85);
	not (d143, d10);
	nor (d144, d93, d108);
	xor (d145, d80, d122);
	nor (d146, d108, d119);
	not (d147, d121);
	buf (d148, d111);
	xor (d149, d99, d106);
	xor (d150, d85, d128);
	xnor (d151, d104, d129);
	not (d152, d126);
	nand (d153, d65, d109);
	nor (d154, d86, d99);
	nand (d155, d67, d79);
	xor (d156, d77, d117);
	or (d157, d76, d127);
	xnor (d158, d71, d114);
	and (d159, d85, d135);
	or (d160, d81, d101);
	not (d161, d94);
	or (d162, d75, d126);
	xnor (d163, d69, d75);
	buf (d164, d30);
	and (d165, d116);
	nor (d166, d72, d114);
	not (d167, d41);
	nor (d168, d80, d112);
	xor (d169, d110, d113);
	nor (d170, d79, d135);
	or (d171, d111, d131);
	buf (d172, d95);
	not (d173, d136);
	or (d174, d87, d130);
	not (d175, d112);
	and (d176, d83, d99);
	or (d177, d71, d82);
	xnor (d178, d91, d119);
	or (d179, d112, d134);
	nand (d180, d83, d108);
	or (d181, d98, d99);
	and (d182, d72, d135);
	buf (d183, d8);
	xor (d184, d75, d111);
	nand (d185, d70, d79);
	nand (d186, d72, d97);
	and (d187, d94, d131);
	nand (d188, d99, d125);
	xnor (d189, d115);
	not (d190, d24);
	xor (d191, d85, d119);
	nor (d192, d114, d116);
	not (d193, d53);
	nand (d194, d88, d90);
	nand (d195, d75, d115);
	not (d196, d2);
	xnor (d197, d107, d114);
	nor (d198, d82, d102);
	xnor (d199, d71, d124);
	buf (d200, d102);
	buf (d201, d100);
	nor (d202, d93, d122);
	nand (d203, d139, d176);
	not (d204, d79);
	or (d205, d175, d185);
	nor (d206, d156, d188);
	buf (d207, d163);
	xor (d208, d159, d167);
	xor (d209, d171, d198);
	or (d210, d192, d201);
	buf (d211, d106);
	nand (d212, d159, d178);
	buf (d213, d48);
	buf (d214, d19);
	xor (d215, d185, d194);
	or (d216, d144, d160);
	nand (d217, d143, d153);
	buf (d218, d162);
	or (d219, d139, d168);
	and (d220, d145, d162);
	and (d221, d167, d182);
	nor (d222, d153, d193);
	not (d223, d191);
	buf (d224, d90);
	xnor (d225, d178, d193);
	and (d226, d142, d146);
	or (d227, d144, d147);
	and (d228, d164, d177);
	not (d229, d76);
	and (d230, d183, d201);
	xor (d231, d138, d187);
	xor (d232, d145, d156);
	nand (d233, d196, d197);
	not (d234, d156);
	buf (d235, d65);
	xnor (d236, d174, d190);
	nor (d237, d150, d172);
	nand (d238, d184, d193);
	xnor (d239, d145, d189);
	xnor (d240, d152, d181);
	nor (d241, d144, d176);
	and (d242, d141, d152);
	xor (d243, d168, d193);
	nand (d244, d173, d196);
	xnor (d245, d143, d185);
	xor (d246, d146, d160);
	xor (d247, d163, d190);
	and (d248, d170, d196);
	nor (d249, d144, d198);
	not (d250, d12);
	xnor (d251, d157, d191);
	buf (d252, d45);
	not (d253, d98);
	nand (d254, d191, d197);
	xor (d255, d217, d224);
	and (d256, d204, d211);
	nor (d257, d224, d226);
	buf (d258, d114);
	xor (d259, d245, d249);
	xnor (d260, d220, d234);
	or (d261, d210, d224);
	nand (d262, d246, d251);
	or (d263, d215, d244);
	or (d264, d218, d250);
	nor (d265, d229, d243);
	not (d266, d159);
	nand (d267, d225, d250);
	xnor (d268, d244, d245);
	or (d269, d213, d244);
	xnor (d270, d211, d249);
	not (d271, d157);
	nor (d272, d215, d254);
	not (d273, d90);
	buf (d274, d68);
	or (d275, d228, d244);
	or (d276, d213, d232);
	nor (d277, d208, d241);
	xor (d278, d229, d233);
	nor (d279, d240, d254);
	xnor (d280, d234, d246);
	xor (d281, d239, d246);
	nor (d282, d241, d242);
	and (d283, d220, d232);
	xor (d284, d210, d244);
	and (d285, d220, d228);
	xor (d286, d230, d238);
	xnor (d287, d214, d233);
	buf (d288, d203);
	xnor (d289, d235, d237);
	and (d290, d227, d251);
	or (d291, d227, d228);
	nor (d292, d222, d229);
	nor (d293, d227, d247);
	and (d294, d208, d236);
	buf (d295, d165);
	nor (d296, d228, d232);
	or (d297, d230, d236);
	nand (d298, d234, d247);
	xnor (d299, d209, d218);
	nand (d300, d206, d252);
	xor (d301, d220, d236);
	or (d302, d216, d253);
	xor (d303, d203, d207);
	or (d304, d222, d224);
	xor (d305, d219, d237);
	buf (d306, d152);
	xor (d307, d203, d206);
	xnor (d308, d217, d231);
	and (d309, d209, d221);
	nor (d310, d235, d237);
	nand (d311, d204, d243);
	nand (d312, d215, d218);
	buf (d313, d40);
	nor (d314, d208, d240);
	nor (d315, d263, d278);
	and (d316, d256, d271);
	and (d317, d281, d288);
	xor (d318, d285, d291);
	not (d319, d241);
	and (d320, d284, d286);
	xor (d321, d260, d305);
	not (d322, d141);
	nor (d323, d303, d308);
	buf (d324, d257);
	and (d325, d297, d313);
	xor (d326, d277, d314);
	and (d327, d299, d301);
	and (d328, d286, d303);
	xnor (d329, d277, d295);
	or (d330, d296, d312);
	nand (d331, d277, d305);
	nand (d332, d283, d303);
	and (d333, d279, d285);
	or (d334, d261, d313);
	nor (d335, d266, d269);
	buf (d336, d37);
	buf (d337, d160);
	buf (d338, d88);
	xnor (d339, d280, d297);
	xor (d340, d285, d302);
	and (d341, d267, d296);
	nor (d342, d306, d313);
	and (d343, d258, d298);
	xnor (d344, d270, d310);
	xnor (d345, d277, d305);
	xor (d346, d259, d262);
	buf (d347, d239);
	or (d348, d299, d308);
	not (d349, d216);
	buf (d350, d126);
	xor (d351, d262, d290);
	xnor (d352, d276, d300);
	or (d353, d267, d280);
	buf (d354, d292);
	xnor (d355, d275, d282);
	nor (d356, d259, d294);
	xor (d357, d271, d280);
	and (d358, d299, d313);
	not (d359, d119);
	nand (d360, d262, d266);
	and (d361, d264, d298);
	not (d362, d294);
	or (d363, d284, d310);
	or (d364, d279, d287);
	and (d365, d259, d314);
	xnor (d366, d280, d296);
	nand (d367, d269, d296);
	xnor (d368, d273, d288);
	nand (d369, d279, d310);
	nand (d370, d269, d312);
	and (d371, d268, d313);
	nor (d372, d258, d278);
	or (d373, d297, d298);
	nor (d374, d267, d299);
	nor (d375, d261, d267);
	or (d376, d274, d286);
	not (d377, d128);
	xor (d378, d286, d287);
	and (d379, d286, d305);
	not (d380, d309);
	or (d381, d263, d292);
	xor (d382, d267, d273);
	xor (d383, d274, d292);
	buf (d384, d262);
	xnor (d385, d328, d377);
	or (d386, d320, d325);
	xor (d387, d318, d372);
	nor (d388, d344, d359);
	and (d389, d347, d351);
	not (d390, d100);
	not (d391, d202);
	nor (d392, d330, d377);
	nand (d393, d330, d377);
	not (d394, d353);
	buf (d395, d3);
	nor (d396, d331, d360);
	xor (d397, d391, d393);
	nand (d398, d387, d395);
	nor (d399, d387, d388);
	buf (d400, d118);
	and (d401, d386);
	xnor (d402, d388, d392);
	nor (d403, d393, d395);
	or (d404, d386, d393);
	not (d405, d149);
	not (d406, d210);
	nor (d407, d385, d389);
	nor (d408, d385, d396);
	xor (d409, d388, d389);
	not (d410, d189);
	xor (d411, d387, d393);
	nor (d412, d385, d386);
	or (d413, d385, d395);
	nor (d414, d389, d394);
	and (d415, d385, d394);
	nand (d416, d389, d394);
	xnor (d417, d389, d393);
	xnor (d418, d390, d391);
	buf (d419, d251);
	nor (d420, d390, d393);
	xor (d421, d389, d390);
	not (d422, d39);
	not (d423, d35);
	buf (d424, d345);
	buf (d425, d171);
	and (d426, d392, d394);
	buf (d427, d129);
	buf (d428, d124);
	nand (d429, d393, d394);
	not (d430, d118);
	and (d431, d391, d395);
	xnor (d432, d395, d396);
	xnor (d433, d387, d396);
	nand (d434, d390, d392);
	buf (d435, d176);
	or (d436, d387, d391);
	or (d437, d389);
	xor (d438, d393, d395);
	nand (d439, d390, d391);
	nand (d440, d393, d395);
	nor (d441, d386, d394);
	or (d442, d385, d391);
	xnor (d443, d393, d394);
	or (d444, d387);
	buf (d445, d204);
	and (d446, d386, d388);
	not (d447, d296);
	not (d448, d80);
	xnor (d449, d387, d394);
	and (d450, d386, d390);
	or (d451, d390, d396);
	nor (d452, d385, d387);
	xnor (d453, d385, d392);
	buf (d454, d339);
	nor (d455, d387, d389);
	xor (d456, d389, d392);
	nand (d457, d424, d445);
	xor (d458, d424, d425);
	or (d459, d400, d422);
	and (d460, d398, d427);
	xnor (d461, d442, d455);
	nand (d462, d418, d456);
	xor (d463, d420, d428);
	and (d464, d403, d439);
	xor (d465, d415, d446);
	nor (d466, d408, d430);
	or (d467, d431, d446);
	xnor (d468, d430, d453);
	or (d469, d410, d442);
	nor (d470, d444, d452);
	xor (d471, d413, d427);
	not (d472, d304);
	nand (d473, d427, d446);
	and (d474, d415, d442);
	nor (d475, d415, d445);
	buf (d476, d375);
	nand (d477, d405, d440);
	not (d478, d50);
	and (d479, d427, d446);
	nor (d480, d435, d438);
	not (d481, d323);
	not (d482, d282);
	and (d483, d404, d421);
	or (d484, d421, d456);
	buf (d485, d244);
	not (d486, d273);
	nand (d487, d414, d448);
	xnor (d488, d407, d454);
	not (d489, d343);
	nand (d490, d409, d428);
	xor (d491, d429, d453);
	not (d492, d104);
	nand (d493, d429, d446);
	and (d494, d429, d447);
	and (d495, d414, d437);
	nand (d496, d430, d437);
	nand (d497, d437, d444);
	not (d498, d198);
	and (d499, d435, d451);
	and (d500, d419, d423);
	and (d501, d405, d446);
	nor (d502, d442, d456);
	nor (d503, d435, d441);
	or (d504, d419, d420);
	and (d505, d414, d416);
	not (d506, d176);
	xor (d507, d412, d427);
	xnor (d508, d398, d447);
	nor (d509, d410, d412);
	xor (d510, d411, d426);
	buf (d511, d404);
	xnor (d512, d410, d439);
	not (d513, d32);
	buf (d514, d93);
	nor (d515, d397, d419);
	xnor (d516, d468, d478);
	and (d517, d459, d485);
	xnor (d518, d462, d503);
	xnor (d519, d473, d502);
	and (d520, d477, d499);
	buf (d521, d376);
	nor (d522, d457, d476);
	not (d523, d288);
	nor (d524, d457, d465);
	nor (d525, d470, d508);
	buf (d526, d369);
	and (d527, d461, d503);
	not (d528, d144);
	xor (d529, d474, d475);
	buf (d530, d446);
	xor (d531, d471, d478);
	or (d532, d474, d512);
	or (d533, d487, d493);
	or (d534, d470, d504);
	nand (d535, d505, d507);
	and (d536, d470, d487);
	xnor (d537, d486, d506);
	xor (d538, d465, d493);
	nand (d539, d482, d503);
	xor (d540, d458, d479);
	nor (d541, d472, d479);
	xor (d542, d459, d497);
	or (d543, d468, d483);
	nor (d544, d474, d477);
	xor (d545, d487, d499);
	buf (d546, d295);
	xnor (d547, d497, d511);
	nor (d548, d486, d515);
	nor (d549, d471, d503);
	buf (d550, d144);
	buf (d551, d258);
	or (d552, d489, d506);
	xnor (d553, d489, d510);
	nor (d554, d470, d497);
	nor (d555, d457, d513);
	nor (d556, d487, d494);
	xor (d557, d461, d504);
	xnor (d558, d459, d472);
	not (d559, d345);
	or (d560, d461, d473);
	or (d561, d461, d496);
	or (d562, d497, d504);
	nor (d563, d468, d474);
	nand (d564, d457, d492);
	xnor (d565, d474, d493);
	not (d566, d221);
	buf (d567, d74);
	xnor (d568, d485, d494);
	nor (d569, d464, d506);
	nand (d570, d462, d501);
	or (d571, d513);
	buf (d572, d300);
	nand (d573, d478, d491);
	nand (d574, d497);
	xor (d575, d465, d503);
	or (d576, d493, d507);
	or (d577, d457, d515);
	buf (d578, d206);
	nand (d579, d497, d500);
	nand (d580, d484, d487);
	xnor (d581, d511);
	xnor (d582, d466, d510);
	nand (d583, d504, d508);
	nand (d584, d468, d498);
	xnor (d585, d470, d492);
	assign f1 = d547;
	assign f2 = d546;
	assign f3 = d528;
	assign f4 = d581;
	assign f5 = d526;
	assign f6 = d524;
	assign f7 = d561;
	assign f8 = d542;
	assign f9 = d545;
	assign f10 = d557;
	assign f11 = d519;
	assign f12 = d526;
endmodule
