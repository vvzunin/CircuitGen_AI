module CCGRCG40( x0, x1, x2, f1, f2, f3 );

	input x0, x1, x2;
	output f1, f2, f3;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263;

	or (d1, x1, x2);
	not (d2, x1);
	nor (d3, x0, x1);
	xnor (d4, x1, x2);
	nand (d5, x0, x1);
	xor (d6, x0, x2);
	not (d7, x0);
	xor (d8, x0);
	or (d9, x1);
	xnor (d10, x0, x2);
	or (d11, x0);
	and (d12, x1);
	buf (d13, x2);
	or (d14, x2);
	and (d15, x0, x1);
	xnor (d16, x0, x1);
	and (d17, x1, x2);
	xor (d18, x0, x1);
	xor (d19, x1, x2);
	xnor (d20, x0, x1);
	xnor (d21, x2);
	or (d22, x0, x2);
	nor (d23, x0);
	buf (d24, x0);
	nand (d25, x2);
	not (d26, x2);
	and (d27, x0);
	xnor (d28, x1, x2);
	nor (d29, x0, x2);
	nand (d30, x0, x1);
	and (d31, x0, x2);
	xnor (d32, x0, x2);
	nor (d33, x1);
	or (d34, d3, d15);
	not (d35, d17);
	xnor (d36, d5, d32);
	xnor (d37, d10, d15);
	xor (d38, d14, d28);
	and (d39, d5, d30);
	and (d40, d10, d11);
	not (d41, d6);
	nand (d42, d4, d26);
	nor (d43, d11, d12);
	xor (d44, d30);
	nand (d45, d1, d8);
	buf (d46, d7);
	nor (d47, d10, d18);
	and (d48, d13, d18);
	nand (d49, d7, d12);
	buf (d50, d12);
	xnor (d51, d10, d26);
	nor (d52, d11, d26);
	or (d53, d2, d30);
	xnor (d54, d13, d31);
	buf (d55, d16);
	and (d56, d24, d32);
	and (d57, d15, d21);
	nor (d58, d8, d17);
	xor (d59, d25, d27);
	xor (d60, d2, d14);
	and (d61, d5, d6);
	not (d62, d16);
	or (d63, d23, d32);
	or (d64, d11, d16);
	or (d65, d22, d28);
	xnor (d66, d4, d33);
	xor (d67, d6, d17);
	and (d68, d30, d33);
	and (d69, d2, d4);
	not (d70, d5);
	nand (d71, d1, d28);
	nor (d72, d10, d29);
	nor (d73, d22, d24);
	xor (d74, d8, d25);
	and (d75, d12, d19);
	nor (d76, d35, d57);
	xnor (d77, d47, d71);
	xnor (d78, d57, d68);
	or (d79, d41, d72);
	xnor (d80, d48, d50);
	not (d81, d74);
	xor (d82, d35, d74);
	or (d83, d46, d49);
	and (d84, d40, d56);
	xnor (d85, d44, d67);
	buf (d86, d28);
	nand (d87, d56, d62);
	and (d88, d38, d52);
	nand (d89, d44, d55);
	xor (d90, d41, d50);
	nand (d91, d34, d55);
	and (d92, d35, d58);
	xor (d93, d64, d66);
	nand (d94, d38, d74);
	nor (d95, d53, d56);
	xnor (d96, d50, d72);
	nor (d97, d48, d74);
	xor (d98, d53, d67);
	xor (d99, d44, d69);
	nor (d100, d61, d65);
	nand (d101, d44, d61);
	xor (d102, d51, d72);
	or (d103, d48, d73);
	and (d104, d68, d74);
	nand (d105, d53, d60);
	xor (d106, d38, d47);
	not (d107, d59);
	nand (d108, d42, d60);
	not (d109, d30);
	not (d110, d55);
	or (d111, d53, d59);
	nand (d112, d61, d68);
	buf (d113, d22);
	xor (d114, d45, d49);
	nor (d115, d35, d62);
	and (d116, d36, d62);
	xor (d117, d63, d74);
	or (d118, d49, d64);
	xor (d119, d37, d69);
	nor (d120, d38, d74);
	not (d121, d27);
	buf (d122, d18);
	and (d123, d100, d109);
	or (d124, d79, d97);
	not (d125, d119);
	not (d126, d41);
	not (d127, d107);
	nor (d128, d89, d111);
	nor (d129, d90, d112);
	and (d130, d109, d118);
	xor (d131, d109, d114);
	or (d132, d84, d89);
	nor (d133, d103, d108);
	or (d134, d90, d102);
	and (d135, d78, d121);
	nand (d136, d102, d119);
	nor (d137, d103, d119);
	nand (d138, d99);
	nand (d139, d96, d121);
	or (d140, d132, d137);
	nand (d141, d134, d137);
	and (d142, d129, d135);
	xor (d143, d131, d137);
	and (d144, d130, d138);
	not (d145, d83);
	nor (d146, d126, d137);
	and (d147, d126, d132);
	nor (d148, d128, d136);
	xor (d149, d128, d129);
	xnor (d150, d127, d129);
	xnor (d151, d128, d134);
	xnor (d152, d123, d139);
	xor (d153, d134, d139);
	not (d154, d34);
	not (d155, d136);
	nand (d156, d135, d138);
	xor (d157, d123, d132);
	nor (d158, d124);
	xnor (d159, d130, d135);
	xor (d160, d123, d125);
	nor (d161, d135, d138);
	or (d162, d124, d133);
	nor (d163, d130, d136);
	xor (d164, d132, d138);
	or (d165, d137, d138);
	nor (d166, d127, d130);
	or (d167, d130, d131);
	nand (d168, d131, d136);
	buf (d169, d1);
	xor (d170, d130, d132);
	or (d171, d126, d131);
	xnor (d172, d125, d135);
	xor (d173, d135, d136);
	and (d174, d125, d127);
	nand (d175, d129, d135);
	nor (d176, d131, d136);
	and (d177, d134, d136);
	xnor (d178, d128, d136);
	buf (d179, d119);
	nor (d180, d123, d124);
	xnor (d181, d131, d139);
	nor (d182, d125, d128);
	xor (d183, d130, d138);
	not (d184, d98);
	or (d185, d140, d172);
	nand (d186, d160, d167);
	and (d187, d144, d157);
	xor (d188, d170, d178);
	nor (d189, d149, d168);
	or (d190, d169, d172);
	buf (d191, d64);
	xnor (d192, d154, d167);
	nand (d193, d143, d165);
	or (d194, d143, d172);
	not (d195, d128);
	buf (d196, d92);
	nand (d197, d170, d179);
	or (d198, d174, d179);
	or (d199, d147, d176);
	buf (d200, d176);
	xor (d201, d164, d172);
	and (d202, d155, d169);
	buf (d203, d48);
	buf (d204, d144);
	nor (d205, d166, d170);
	nand (d206, d157, d180);
	or (d207, d145, d153);
	nand (d208, d142, d176);
	not (d209, d167);
	xnor (d210, d148, d158);
	xor (d211, d161, d173);
	nand (d212, d149, d171);
	nor (d213, d168, d176);
	and (d214, d146, d153);
	not (d215, d78);
	nand (d216, d175, d182);
	nor (d217, d168, d183);
	and (d218, d145, d175);
	xor (d219, d151, d166);
	nor (d220, d147, d177);
	xor (d221, d164, d176);
	xor (d222, d142, d158);
	xor (d223, d160, d181);
	xnor (d224, d150, d178);
	or (d225, d170, d181);
	xnor (d226, d155, d162);
	xnor (d227, d150, d164);
	and (d228, d147, d150);
	nand (d229, d170, d180);
	nand (d230, d140, d149);
	xor (d231, d148, d153);
	and (d232, d151, d181);
	nand (d233, d145, d147);
	or (d234, d150, d158);
	nor (d235, d149, d155);
	xnor (d236, d164);
	or (d237, d142, d151);
	buf (d238, d96);
	or (d239, d153, d175);
	xor (d240, d149, d175);
	nor (d241, d157, d159);
	xor (d242, d150, d172);
	and (d243, d143, d176);
	xor (d244, d178, d181);
	buf (d245, d26);
	xor (d246, d140, d166);
	or (d247, d141, d169);
	xnor (d248, d158, d183);
	xnor (d249, d142, d143);
	xnor (d250, d153, d162);
	or (d251, d170, d172);
	nor (d252, d143, d168);
	xor (d253, d142, d162);
	or (d254, d154, d172);
	xnor (d255, d147, d171);
	xnor (d256, d143, d155);
	xnor (d257, d164, d183);
	nand (d258, d173, d179);
	nand (d259, d157, d178);
	not (d260, d114);
	xor (d261, d152, d163);
	not (d262, d88);
	buf (d263, d82);
	assign f1 = d188;
	assign f2 = d194;
	assign f3 = d213;
endmodule
