module CCGRCG194( x0, x1, x2, x3, x4, x5, x6, f1, f2, f3, f4 );

	input x0, x1, x2, x3, x4, x5, x6;
	output f1, f2, f3, f4;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209;

	nand (d1, x2, x3);
	nand (d2, x1, x3);
	nand (d3, x1, x6);
	xnor (d4, x5, x6);
	not (d5, x1);
	or (d6, x4, x5);
	and (d7, x1, x6);
	or (d8, x3, x5);
	buf (d9, x5);
	xnor (d10, x2);
	or (d11, x3, x6);
	and (d12, x1, x3);
	xor (d13, x3, x5);
	nand (d14, x5);
	nand (d15, x3, x5);
	or (d16, x1, x6);
	nand (d17, x1);
	and (d18, x1, x5);
	nand (d19, x1, x3);
	or (d20, x3, x4);
	nand (d21, x0, x4);
	not (d22, x3);
	xor (d23, x3, x4);
	xor (d24, x1, x6);
	xor (d25, x0, x3);
	not (d26, x2);
	and (d27, x5, x6);
	nor (d28, x0, x2);
	or (d29, x4, x5);
	xnor (d30, x2, x5);
	xor (d31, x1, x5);
	nor (d32, x2, x6);
	nand (d33, x4);
	nor (d34, x5);
	xor (d35, x1, x4);
	or (d36, x2);
	nor (d37, x4, x5);
	not (d38, x5);
	nand (d39, x0, x2);
	or (d40, x1, x2);
	nor (d41, x3, x6);
	and (d42, x1, x2);
	buf (d43, x4);
	or (d44, x2, x6);
	xnor (d45, x1, x2);
	not (d46, x0);
	xnor (d47, x1, x3);
	xor (d48, x1, x5);
	buf (d49, x3);
	or (d50, x1, x4);
	nand (d51, x1, x4);
	nand (d52, x3, x6);
	nor (d53, x2, x5);
	not (d54, x6);
	xnor (d55, x3);
	or (d56, x0, x2);
	xor (d57, x0, x4);
	nor (d58, x0, x4);
	xor (d59, x3, x6);
	buf (d60, x0);
	buf (d61, x1);
	and (d62, x0, x3);
	or (d63, x0, x5);
	nor (d64, d4, d9);
	nor (d65, d36, d43);
	xor (d66, d4, d33);
	xor (d67, d19, d47);
	xor (d68, d36, d62);
	xnor (d69, d44, d50);
	or (d70, d10, d38);
	nor (d71, d2, d14);
	xor (d72, d5, d42);
	nor (d73, d32, d52);
	xnor (d74, d11, d38);
	xor (d75, d3, d58);
	or (d76, d24, d61);
	buf (d77, x2);
	xor (d78, d38, d39);
	or (d79, d25, d38);
	not (d80, d6);
	and (d81, d41, d50);
	nor (d82, d66, d74);
	xor (d83, d79, d81);
	xnor (d84, d72, d80);
	xor (d85, d70, d74);
	xor (d86, d69, d79);
	xor (d87, d65, d77);
	nor (d88, d64, d77);
	or (d89, d71, d81);
	nand (d90, d75, d78);
	and (d91, d78, d80);
	xor (d92, d67, d79);
	buf (d93, d23);
	and (d94, d71, d80);
	xor (d95, d69, d79);
	xnor (d96, d70, d74);
	nor (d97, d64, d69);
	buf (d98, d11);
	not (d99, d31);
	xor (d100, d71, d74);
	nand (d101, d64, d68);
	and (d102, d67, d71);
	not (d103, d72);
	or (d104, d69, d73);
	buf (d105, d80);
	nand (d106, d73, d78);
	xnor (d107, d69, d71);
	and (d108, d72, d81);
	not (d109, d32);
	not (d110, d75);
	or (d111, d70, d79);
	nand (d112, d72, d80);
	buf (d113, d70);
	and (d114, d71, d80);
	xnor (d115, d77, d79);
	nand (d116, d70, d78);
	or (d117, d65, d74);
	or (d118, d64, d67);
	and (d119, d76, d78);
	nor (d120, d73, d78);
	xor (d121, d67, d75);
	xnor (d122, d71, d80);
	not (d123, d79);
	or (d124, d64, d81);
	nor (d125, d75, d77);
	and (d126, d71, d75);
	nor (d127, d73, d74);
	nor (d128, d76);
	buf (d129, d5);
	buf (d130, d41);
	or (d131, d67, d76);
	xnor (d132, d76, d80);
	and (d133, d90, d132);
	and (d134, d100, d112);
	nor (d135, d84, d92);
	or (d136, d85, d123);
	xnor (d137, d99, d129);
	nor (d138, d114, d122);
	not (d139, d20);
	and (d140, d139);
	or (d141, d133, d139);
	nor (d142, d135);
	nor (d143, d135, d138);
	and (d144, d137);
	and (d145, d135, d138);
	nor (d146, d133, d137);
	buf (d147, d121);
	or (d148, d133, d137);
	buf (d149, d45);
	or (d150, d135);
	not (d151, d35);
	xnor (d152, d133, d138);
	not (d153, d65);
	xor (d154, d135, d137);
	nor (d155, d133, d136);
	and (d156, d138, d139);
	buf (d157, d42);
	nor (d158, d137, d138);
	nand (d159, d134, d139);
	buf (d160, d73);
	nor (d161, d134, d135);
	nor (d162, d141, d145);
	buf (d163, d127);
	xnor (d164, d145, d159);
	buf (d165, d48);
	xor (d166, d143);
	not (d167, d137);
	buf (d168, d123);
	not (d169, d38);
	not (d170, d73);
	nand (d171, d145, d152);
	not (d172, d148);
	xnor (d173, d142, d158);
	or (d174, d144, d151);
	nand (d175, d143, d160);
	or (d176, d159);
	buf (d177, d69);
	not (d178, d96);
	and (d179, d168, d177);
	nor (d180, d169, d178);
	nor (d181, d162, d176);
	xor (d182, d168, d169);
	and (d183, d166, d173);
	and (d184, d174, d178);
	or (d185, d166, d169);
	nand (d186, d169, d171);
	xnor (d187, d174, d175);
	nand (d188, d169, d172);
	or (d189, d163, d170);
	nor (d190, d164, d178);
	nor (d191, d162, d171);
	nand (d192, d187, d190);
	and (d193, d180, d184);
	or (d194, d180);
	xnor (d195, d185, d187);
	xnor (d196, d180, d191);
	buf (d197, d2);
	nor (d198, d180, d184);
	buf (d199, d166);
	and (d200, d179, d188);
	nor (d201, d181, d190);
	xor (d202, d179, d183);
	nor (d203, d179, d185);
	or (d204, d180, d182);
	and (d205, d180, d182);
	xor (d206, d187, d189);
	xor (d207, d180, d185);
	nor (d208, d180, d188);
	xor (d209, d179, d180);
	assign f1 = d200;
	assign f2 = d209;
	assign f3 = d208;
	assign f4 = d197;
endmodule
