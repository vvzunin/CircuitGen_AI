module CCGRCG31( x0, x1, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17 );

	input x0, x1;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201;

	or (d1, x0);
	xor (d2, x0, x1);
	and (d3, x0, x1);
	nand (d4, x1);
	xor (d5, x0);
	nor (d6, x1);
	xor (d7, x0, x1);
	not (d8, x0);
	nor (d9, x0, x1);
	buf (d10, x0);
	and (d11, x0, x1);
	or (d12, x0, x1);
	xnor (d13, x0, x1);
	buf (d14, x1);
	nor (d15, d1, d7);
	buf (d16, d9);
	or (d17, d7, d8);
	xnor (d18, d7, d11);
	buf (d19, d11);
	buf (d20, d12);
	xor (d21, d1, d3);
	nand (d22, d13);
	nor (d23, d1, d14);
	not (d24, d3);
	not (d25, d11);
	not (d26, d13);
	xnor (d27, d4, d9);
	and (d28, d9, d13);
	nand (d29, d6, d10);
	and (d30, d9);
	and (d31, d3, d11);
	or (d32, d13, d14);
	xor (d33, d10, d12);
	nand (d34, d1, d9);
	and (d35, d2, d4);
	or (d36, d2, d13);
	xnor (d37, d17, d26);
	nand (d38, d16, d25);
	nor (d39, d18, d31);
	nand (d40, d20, d33);
	xor (d41, d17, d26);
	buf (d42, d20);
	xnor (d43, d20, d23);
	nor (d44, d18, d28);
	and (d45, d16, d28);
	xor (d46, d20, d36);
	xor (d47, d23, d34);
	not (d48, d35);
	xor (d49, d25, d27);
	nand (d50, d18, d23);
	and (d51, d15, d30);
	nor (d52, d21, d22);
	xor (d53, d18, d21);
	nor (d54, d29, d31);
	or (d55, d19, d26);
	and (d56, d25);
	and (d57, d18, d23);
	xnor (d58, d16, d19);
	buf (d59, d29);
	not (d60, d20);
	xnor (d61, d23, d26);
	nor (d62, d34);
	nand (d63, d28, d30);
	not (d64, d10);
	or (d65, d15, d30);
	not (d66, d34);
	and (d67, d18, d29);
	nor (d68, d16, d24);
	xor (d69, d21, d23);
	and (d70, d32, d36);
	xor (d71, d19, d26);
	nor (d72, d25, d34);
	xor (d73, d22, d31);
	nor (d74, d24, d35);
	buf (d75, d3);
	and (d76, d34, d36);
	nor (d77, d17, d28);
	nor (d78, d18, d24);
	nor (d79, d16, d27);
	nor (d80, d24, d35);
	not (d81, x1);
	nand (d82, d20, d22);
	or (d83, d19, d22);
	nor (d84, d15, d28);
	and (d85, d20, d21);
	nand (d86, d26, d29);
	and (d87, d19, d34);
	nand (d88, d25, d31);
	nand (d89, d30, d35);
	nor (d90, d18, d31);
	or (d91, d28, d31);
	xor (d92, d25, d26);
	and (d93, d22, d24);
	nand (d94, d19, d32);
	or (d95, d31, d34);
	nor (d96, d25, d31);
	buf (d97, d1);
	not (d98, d18);
	xor (d99, d33, d36);
	nand (d100, d19, d36);
	nor (d101, d21, d34);
	nand (d102, d58, d71);
	nor (d103, d49, d60);
	xor (d104, d43, d82);
	not (d105, d96);
	or (d106, d76, d101);
	or (d107, d94, d97);
	and (d108, d58, d78);
	buf (d109, d65);
	xnor (d110, d74, d88);
	xor (d111, d105, d109);
	and (d112, d107);
	and (d113, d102, d106);
	xor (d114, d103, d108);
	and (d115, d108);
	xor (d116, d109);
	xnor (d117, d108, d109);
	xor (d118, d103, d105);
	not (d119, d38);
	or (d120, d103, d110);
	nand (d121, d108);
	nor (d122, d104, d110);
	buf (d123, d70);
	xnor (d124, d108, d109);
	or (d125, d110);
	and (d126, d102, d104);
	xor (d127, d107);
	nor (d128, d106, d109);
	xor (d129, d104, d106);
	buf (d130, d17);
	xor (d131, d105, d110);
	nor (d132, d102, d109);
	nor (d133, d102, d105);
	not (d134, d57);
	or (d135, d107);
	or (d136, d102, d103);
	and (d137, d103, d110);
	nand (d138, d103, d108);
	and (d139, d109);
	xnor (d140, d102, d110);
	xor (d141, d105, d110);
	buf (d142, d33);
	buf (d143, d73);
	or (d144, d102, d107);
	nor (d145, d104, d105);
	or (d146, d105, d109);
	not (d147, d61);
	xnor (d148, d107, d108);
	and (d149, d105, d107);
	xnor (d150, d102, d105);
	or (d151, d104);
	not (d152, d43);
	nand (d153, d107, d109);
	nor (d154, d105, d109);
	and (d155, d106, d110);
	xnor (d156, d102, d104);
	buf (d157, d54);
	not (d158, d88);
	xnor (d159, d103, d110);
	xnor (d160, d102, d107);
	nor (d161, d105, d110);
	xor (d162, d102, d105);
	or (d163, d103, d104);
	not (d164, d53);
	xnor (d165, d104, d108);
	xnor (d166, d106, d110);
	xnor (d167, d103, d106);
	buf (d168, d44);
	xnor (d169, d109);
	xor (d170, d105, d109);
	xnor (d171, d103, d104);
	nand (d172, d104, d108);
	nand (d173, d104, d105);
	not (d174, d73);
	nor (d175, d102, d108);
	or (d176, d107, d109);
	not (d177, d80);
	nor (d178, d104, d107);
	and (d179, d103, d106);
	nand (d180, d103, d106);
	nor (d181, d102, d108);
	xor (d182, d103, d108);
	not (d183, d85);
	not (d184, d50);
	and (d185, d108, d109);
	nand (d186, d103, d109);
	xnor (d187, d102);
	nor (d188, d104, d108);
	nand (d189, d105);
	and (d190, d102, d104);
	buf (d191, d62);
	xnor (d192, d107, d109);
	nand (d193, d104);
	and (d194, d108, d109);
	nor (d195, d105, d108);
	xnor (d196, d103, d105);
	xor (d197, d103, d104);
	or (d198, d102, d107);
	and (d199, d106, d107);
	nand (d200, d103, d108);
	xor (d201, d107, d108);
	assign f1 = d165;
	assign f2 = d156;
	assign f3 = d167;
	assign f4 = d121;
	assign f5 = d157;
	assign f6 = d181;
	assign f7 = d137;
	assign f8 = d191;
	assign f9 = d179;
	assign f10 = d113;
	assign f11 = d113;
	assign f12 = d189;
	assign f13 = d114;
	assign f14 = d140;
	assign f15 = d158;
	assign f16 = d183;
	assign f17 = d197;
endmodule
