module CCGRCG66( x0, x1, x2, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16 );

	input x0, x1, x2;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314, d315, d316, d317, d318, d319, d320, d321, d322, d323, d324, d325, d326, d327, d328, d329, d330, d331, d332, d333;

	xnor (d1, x1, x2);
	nand (d2, x1, x2);
	or (d3, x0, x2);
	buf (d4, x1);
	nand (d5, x1, x2);
	and (d6, x0, x2);
	and (d7, x0, x1);
	or (d8, x1, x2);
	not (d9, x0);
	not (d10, x2);
	and (d11, x1);
	or (d12, x2);
	nor (d13, x1, x2);
	xnor (d14, x0, x1);
	buf (d15, x2);
	or (d16, x0, x2);
	or (d17, x0, x1);
	not (d18, x1);
	nand (d19, x0);
	xnor (d20, x1, x2);
	buf (d21, x0);
	and (d22, x2);
	or (d23, x0);
	and (d24, x1, x2);
	nand (d25, x2);
	or (d26, x1, x2);
	xor (d27, x1, x2);
	nor (d28, x1);
	xnor (d29, d3, d9);
	xor (d30, d13, d20);
	and (d31, d19, d22);
	not (d32, d14);
	nor (d33, d10, d17);
	xor (d34, d19, d23);
	nand (d35, d18, d20);
	nor (d36, d10, d17);
	xor (d37, d2, d3);
	not (d38, d10);
	xor (d39, d11, d21);
	xor (d40, d3, d6);
	xnor (d41, d10, d21);
	not (d42, d17);
	buf (d43, d4);
	nor (d44, d12, d23);
	nand (d45, d4, d19);
	buf (d46, d28);
	not (d47, d15);
	xnor (d48, d22, d25);
	not (d49, d26);
	xnor (d50, d3, d10);
	xnor (d51, d2, d13);
	xnor (d52, d6, d22);
	xnor (d53, d25, d28);
	buf (d54, d25);
	xnor (d55, d7, d10);
	or (d56, d12, d20);
	and (d57, d7, d27);
	buf (d58, d24);
	or (d59, d12, d21);
	xor (d60, d8, d19);
	and (d61, d13, d28);
	nor (d62, d12, d16);
	xnor (d63, d10, d23);
	nand (d64, d14, d21);
	nand (d65, d12, d23);
	xor (d66, d1, d3);
	nor (d67, d1, d18);
	nor (d68, d14, d19);
	xnor (d69, d2, d27);
	xor (d70, d8, d16);
	and (d71, d19, d27);
	or (d72, d1, d4);
	nor (d73, d14);
	nand (d74, d4, d22);
	or (d75, d13, d23);
	nand (d76, d22, d23);
	xnor (d77, d14, d26);
	and (d78, d9, d15);
	xor (d79, d4, d23);
	xnor (d80, d8, d20);
	or (d81, d10, d14);
	xnor (d82, d3, d20);
	xnor (d83, d8, d9);
	xor (d84, d18, d28);
	not (d85, d16);
	xor (d86, d35, d83);
	nand (d87, d37, d81);
	not (d88, d1);
	and (d89, d52, d58);
	or (d90, d29, d31);
	or (d91, d61, d70);
	and (d92, d31, d47);
	nand (d93, d54, d72);
	not (d94, d33);
	buf (d95, d72);
	buf (d96, d40);
	nor (d97, d43, d74);
	xor (d98, d36, d85);
	nand (d99, d32, d80);
	nand (d100, d56, d78);
	and (d101, d43, d57);
	xor (d102, d34, d51);
	or (d103, d60, d65);
	buf (d104, d34);
	xnor (d105, d47, d84);
	xnor (d106, d78, d84);
	xnor (d107, d63, d73);
	buf (d108, d6);
	nor (d109, d29, d38);
	buf (d110, d10);
	or (d111, d34, d77);
	xor (d112, d47, d85);
	nor (d113, d36, d84);
	nand (d114, d52, d54);
	xnor (d115, d51, d67);
	or (d116, d74, d84);
	buf (d117, d43);
	xnor (d118, d35, d36);
	nand (d119, d33, d47);
	not (d120, d65);
	xnor (d121, d31, d84);
	or (d122, d52, d71);
	nor (d123, d44, d85);
	buf (d124, d80);
	not (d125, d35);
	xnor (d126, d34, d38);
	nor (d127, d54, d68);
	or (d128, d47, d67);
	buf (d129, d29);
	nand (d130, d61, d69);
	or (d131, d44, d64);
	or (d132, d51, d74);
	xor (d133, d42, d59);
	xor (d134, d40);
	not (d135, d2);
	and (d136, d37, d51);
	nor (d137, d42, d75);
	nor (d138, d75, d83);
	not (d139, d79);
	nand (d140, d33, d74);
	and (d141, d70, d75);
	and (d142, d38, d75);
	or (d143, d55, d64);
	or (d144, d32, d56);
	xnor (d145, d34, d57);
	nand (d146, d47, d54);
	and (d147, d41, d52);
	not (d148, d72);
	xnor (d149, d50, d62);
	nand (d150, d34, d38);
	nand (d151, d40, d60);
	and (d152, d57, d69);
	nand (d153, d47, d62);
	not (d154, d28);
	not (d155, d49);
	nor (d156, d37, d54);
	buf (d157, d37);
	nand (d158, d41, d52);
	and (d159, d78, d82);
	nor (d160, d31, d50);
	and (d161, d51, d80);
	xnor (d162, d64, d84);
	and (d163, d71, d73);
	or (d164, d52, d53);
	xnor (d165, d73, d80);
	xor (d166, d44, d66);
	xnor (d167, d67, d70);
	buf (d168, d69);
	or (d169, d71, d77);
	xnor (d170, d48, d52);
	not (d171, d9);
	nand (d172, d31, d33);
	xnor (d173, d32, d77);
	xor (d174, d40, d42);
	nand (d175, d29, d85);
	or (d176, d79, d81);
	and (d177, d41, d83);
	nand (d178, d87, d156);
	not (d179, d43);
	xor (d180, d119, d152);
	xor (d181, d117, d173);
	xor (d182, d88, d121);
	or (d183, d92, d112);
	xnor (d184, d145, d174);
	nand (d185, d101, d175);
	nor (d186, d92, d123);
	and (d187, d143, d168);
	nand (d188, d87, d88);
	not (d189, d58);
	and (d190, d136, d159);
	and (d191, d137, d139);
	not (d192, d127);
	and (d193, d118, d144);
	nand (d194, d86, d139);
	nand (d195, d95, d117);
	nor (d196, d103, d172);
	or (d197, d100, d171);
	not (d198, d151);
	xor (d199, d113, d117);
	xor (d200, d126, d148);
	not (d201, d96);
	xnor (d202, d110, d131);
	or (d203, d124, d129);
	xnor (d204, d100, d123);
	nor (d205, d106, d169);
	xnor (d206, d143, d164);
	and (d207, d96, d162);
	not (d208, d77);
	nand (d209, d158, d170);
	buf (d210, d18);
	or (d211, d116, d170);
	xnor (d212, d101, d145);
	nor (d213, d105, d173);
	xor (d214, d93, d124);
	xor (d215, d98, d108);
	or (d216, d125, d151);
	nor (d217, d139, d143);
	buf (d218, d116);
	nand (d219, d88, d103);
	and (d220, d105, d154);
	buf (d221, d106);
	or (d222, d102, d165);
	nor (d223, d140, d148);
	buf (d224, d167);
	xor (d225, d205, d220);
	xnor (d226, d220, d223);
	nor (d227, d201, d224);
	buf (d228, d36);
	xor (d229, d187, d221);
	xnor (d230, d199, d224);
	nor (d231, d204, d221);
	not (d232, d191);
	xor (d233, d197, d220);
	and (d234, d188, d219);
	and (d235, d180, d215);
	not (d236, d87);
	xnor (d237, d178, d221);
	nor (d238, d191, d208);
	or (d239, d211, d212);
	and (d240, d211, d218);
	or (d241, d191, d214);
	and (d242, d183, d209);
	and (d243, d182, d192);
	nor (d244, d195, d201);
	not (d245, d123);
	xor (d246, d204, d211);
	buf (d247, d215);
	nor (d248, d197, d205);
	nor (d249, d207);
	buf (d250, d22);
	buf (d251, d193);
	not (d252, d114);
	buf (d253, d157);
	not (d254, d45);
	nor (d255, d187, d218);
	or (d256, d183, d185);
	and (d257, d213, d222);
	nor (d258, d205, d214);
	nand (d259, d179, d212);
	buf (d260, d168);
	nand (d261, d197, d222);
	xor (d262, d189, d199);
	and (d263, d182, d185);
	nor (d264, d207, d219);
	xor (d265, d195, d214);
	not (d266, d152);
	nand (d267, d205, d216);
	xnor (d268, d203, d206);
	nand (d269, d195, d217);
	xnor (d270, d206, d216);
	buf (d271, d136);
	nand (d272, d213, d222);
	buf (d273, d84);
	nor (d274, d212, d222);
	xnor (d275, d191, d192);
	xnor (d276, d183, d221);
	nand (d277, d195, d216);
	nand (d278, d194, d220);
	xnor (d279, d193, d222);
	nor (d280, d192, d208);
	not (d281, d20);
	nor (d282, d187, d199);
	xor (d283, d195, d213);
	and (d284, d200, d218);
	buf (d285, d276);
	not (d286, d150);
	not (d287, d209);
	or (d288, d246, d276);
	nand (d289, d241, d284);
	not (d290, d134);
	buf (d291, d166);
	nor (d292, d232, d269);
	not (d293, d36);
	nor (d294, d233, d255);
	not (d295, d279);
	nand (d296, d239, d255);
	and (d297, d245, d277);
	xnor (d298, d240, d281);
	xnor (d299, d229, d236);
	buf (d300, d253);
	xnor (d301, d260);
	not (d302, d94);
	or (d303, d239, d269);
	not (d304, d144);
	xnor (d305, d265, d266);
	not (d306, d159);
	nand (d307, d237, d251);
	and (d308, d228, d241);
	or (d309, d273, d277);
	nand (d310, d230, d253);
	nor (d311, d235, d269);
	buf (d312, d219);
	nor (d313, d239, d283);
	not (d314, d44);
	buf (d315, d172);
	and (d316, d229, d252);
	nand (d317, d225, d242);
	not (d318, d132);
	and (d319, d255, d272);
	buf (d320, d20);
	nand (d321, d264, d272);
	nand (d322, d225, d239);
	xnor (d323, d231, d272);
	nor (d324, d274, d279);
	xor (d325, d238, d273);
	nor (d326, d264, d280);
	xor (d327, d237, d263);
	xor (d328, d252, d279);
	xor (d329, d277, d283);
	buf (d330, d244);
	or (d331, d256, d279);
	nor (d332, d243, d252);
	not (d333, d206);
	assign f1 = d285;
	assign f2 = d322;
	assign f3 = d333;
	assign f4 = d291;
	assign f5 = d328;
	assign f6 = d328;
	assign f7 = d293;
	assign f8 = d313;
	assign f9 = d295;
	assign f10 = d287;
	assign f11 = d320;
	assign f12 = d310;
	assign f13 = d302;
	assign f14 = d286;
	assign f15 = d326;
	assign f16 = d299;
endmodule
