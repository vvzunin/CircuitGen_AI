module CCGRCG146( x0, x1, x2, x3, x4, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17, f18 );

	input x0, x1, x2, x3, x4;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17, f18;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314, d315, d316, d317, d318, d319, d320, d321, d322, d323, d324, d325, d326, d327, d328, d329, d330, d331, d332, d333, d334, d335, d336, d337, d338, d339, d340, d341, d342, d343, d344, d345, d346, d347, d348, d349, d350, d351, d352, d353, d354, d355, d356, d357, d358, d359, d360, d361, d362, d363, d364, d365, d366, d367, d368, d369, d370, d371, d372, d373, d374, d375, d376, d377, d378, d379, d380, d381, d382, d383, d384, d385, d386, d387, d388, d389, d390, d391, d392, d393, d394, d395, d396, d397, d398, d399, d400, d401;

	nand (d1, x2, x3);
	nor (d2, x1, x3);
	buf (d3, x2);
	nor (d4, x4);
	or (d5, x1, x2);
	nor (d6, x2, x3);
	nand (d7, x2, x3);
	or (d8, x0, x1);
	nand (d9, x4);
	not (d10, x1);
	xnor (d11, x1, x2);
	nand (d12, x0, x3);
	not (d13, x0);
	not (d14, x3);
	and (d15, x1, x2);
	nor (d16, x0, x1);
	and (d17, x3, x4);
	xor (d18, x1);
	and (d19, x0, x2);
	and (d20, x1, x4);
	not (d21, x4);
	not (d22, x2);
	nor (d23, x3, x4);
	or (d24, x0);
	nor (d25, x0, x2);
	or (d26, x1, x2);
	and (d27, x2, x4);
	and (d28, d23, d26);
	xnor (d29, d8, d19);
	xor (d30, d6, d12);
	nor (d31, d8);
	nand (d32, d17, d21);
	nand (d33, d5, d19);
	buf (d34, x4);
	xor (d35, d24, d26);
	buf (d36, d27);
	nor (d37, d1, d24);
	nor (d38, d3, d26);
	and (d39, d12, d27);
	buf (d40, d10);
	and (d41, d1, d16);
	xnor (d42, d13, d23);
	xnor (d43, d10, d24);
	or (d44, d7, d9);
	nor (d45, d2, d16);
	nand (d46, d6, d8);
	nand (d47, d19, d25);
	xnor (d48, d13, d22);
	and (d49, d17, d23);
	xnor (d50, d14, d16);
	or (d51, d32, d50);
	xor (d52, d43, d45);
	or (d53, d37, d38);
	nand (d54, d31, d44);
	nor (d55, d44, d46);
	xnor (d56, d29, d41);
	nor (d57, d33, d38);
	xor (d58, d42, d43);
	not (d59, d8);
	not (d60, d13);
	nand (d61, d39, d50);
	buf (d62, d24);
	xor (d63, d31, d41);
	xor (d64, d35, d50);
	xnor (d65, d44, d45);
	nor (d66, d33, d44);
	nand (d67, d32, d48);
	buf (d68, d15);
	or (d69, d46, d50);
	buf (d70, d46);
	or (d71, d37, d45);
	not (d72, d17);
	not (d73, d43);
	xnor (d74, d28, d45);
	not (d75, d16);
	not (d76, d1);
	buf (d77, d42);
	nor (d78, d36, d45);
	and (d79, d30, d39);
	nor (d80, d29, d43);
	or (d81, d32, d33);
	or (d82, d29, d46);
	nor (d83, d40, d44);
	nor (d84, d28, d37);
	xnor (d85, d42, d46);
	nor (d86, d28, d46);
	nand (d87, d37, d40);
	xor (d88, d40, d50);
	xor (d89, d35, d46);
	xor (d90, d42, d45);
	and (d91, d42, d44);
	buf (d92, d5);
	xor (d93, d30, d41);
	and (d94, d33, d48);
	nor (d95, d34, d47);
	nor (d96, d30, d37);
	xor (d97, d31, d40);
	nor (d98, d32, d37);
	not (d99, d11);
	or (d100, d66, d90);
	not (d101, d81);
	xnor (d102, d82, d96);
	nand (d103, d57, d61);
	xnor (d104, d89, d94);
	nand (d105, d61, d85);
	buf (d106, d86);
	xnor (d107, d65, d95);
	nor (d108, d61, d73);
	buf (d109, d7);
	xor (d110, d72, d97);
	xor (d111, d67, d96);
	not (d112, d61);
	nor (d113, d56, d92);
	buf (d114, d58);
	buf (d115, d19);
	buf (d116, d38);
	nor (d117, d58, d83);
	and (d118, d52, d82);
	nor (d119, d57, d73);
	nor (d120, d71, d78);
	not (d121, d97);
	not (d122, d95);
	or (d123, d64, d72);
	or (d124, d78, d88);
	xnor (d125, d58, d77);
	xor (d126, d55, d61);
	xor (d127, d65, d68);
	nand (d128, d65, d82);
	not (d129, d85);
	or (d130, d57, d75);
	or (d131, d56, d87);
	xor (d132, d70, d80);
	nand (d133, d92, d98);
	and (d134, d53, d98);
	or (d135, d62, d74);
	xor (d136, d56, d61);
	buf (d137, d75);
	xnor (d138, d64, d71);
	xnor (d139, d76, d85);
	xnor (d140, d63, d67);
	and (d141, d76, d87);
	buf (d142, d26);
	xnor (d143, d93, d94);
	and (d144, d51, d92);
	nor (d145, d68, d89);
	nand (d146, d91, d96);
	or (d147, d62, d96);
	and (d148, d69, d97);
	or (d149, d60, d97);
	nor (d150, d77, d79);
	nand (d151, d62, d63);
	xnor (d152, d72, d98);
	buf (d153, d17);
	nor (d154, d87, d94);
	nor (d155, d75, d86);
	buf (d156, d29);
	not (d157, d50);
	not (d158, d79);
	and (d159, d52, d93);
	and (d160, d124, d125);
	buf (d161, d137);
	and (d162, d140, d153);
	or (d163, d101, d138);
	or (d164, d100, d104);
	buf (d165, d139);
	not (d166, d23);
	nor (d167, d117, d120);
	not (d168, d148);
	nand (d169, d104, d156);
	and (d170, d105, d119);
	xnor (d171, d111, d112);
	nor (d172, d141, d149);
	xor (d173, d103, d123);
	and (d174, d124, d126);
	xor (d175, d128, d142);
	not (d176, d105);
	and (d177, d127, d149);
	buf (d178, d52);
	and (d179, d104, d114);
	and (d180, d146, d148);
	nor (d181, d114, d122);
	buf (d182, d45);
	xor (d183, d134, d153);
	xnor (d184, d108, d109);
	buf (d185, d3);
	and (d186, d110, d117);
	nand (d187, d106, d148);
	and (d188, d175, d183);
	nand (d189, d178, d184);
	nand (d190, d173, d177);
	nor (d191, d160, d180);
	xnor (d192, d160, d177);
	nand (d193, d166, d171);
	nand (d194, d163, d171);
	xnor (d195, d179, d180);
	xnor (d196, d174, d182);
	nand (d197, d177, d187);
	and (d198, d166, d187);
	xor (d199, d177, d187);
	nand (d200, d164, d169);
	not (d201, d36);
	or (d202, d174, d180);
	nand (d203, d183, d186);
	buf (d204, x1);
	buf (d205, d152);
	xnor (d206, d179, d184);
	not (d207, d47);
	or (d208, d167, d178);
	xnor (d209, d171, d180);
	and (d210, d169, d179);
	or (d211, d180, d186);
	xnor (d212, d169, d172);
	or (d213, d161, d170);
	xnor (d214, d162, d172);
	not (d215, d161);
	or (d216, d180, d185);
	not (d217, d113);
	xnor (d218, d172, d175);
	not (d219, d126);
	not (d220, d135);
	or (d221, d182, d185);
	xor (d222, d171, d172);
	and (d223, d166, d173);
	nand (d224, d164, d165);
	nand (d225, d173, d186);
	or (d226, d163, d177);
	xnor (d227, d168, d178);
	nor (d228, d180, d182);
	nand (d229, d161, d175);
	and (d230, d170, d174);
	and (d231, d162, d174);
	xor (d232, d169, d173);
	xor (d233, d178, d182);
	nand (d234, d163, d187);
	and (d235, d165, d180);
	nor (d236, d179, d183);
	buf (d237, d182);
	nand (d238, d171, d174);
	xor (d239, d166, d179);
	xnor (d240, d169, d173);
	xor (d241, d161, d174);
	nor (d242, d173, d184);
	xor (d243, d161, d177);
	or (d244, d168, d178);
	and (d245, d167, d179);
	or (d246, d169, d185);
	nor (d247, d183, d187);
	or (d248, d163, d180);
	or (d249, d165, d186);
	or (d250, d164, d172);
	nand (d251, d161, d171);
	nand (d252, d174, d183);
	xnor (d253, d163, d186);
	xnor (d254, d168, d183);
	and (d255, d167, d171);
	or (d256, d160, d171);
	and (d257, d166, d172);
	and (d258, d177, d183);
	not (d259, d172);
	nor (d260, d166, d171);
	not (d261, d10);
	xor (d262, d163, d177);
	xnor (d263, d170, d175);
	and (d264, d183, d185);
	or (d265, d165, d169);
	not (d266, d12);
	buf (d267, d16);
	xnor (d268, d162, d171);
	xnor (d269, d178);
	or (d270, d161, d179);
	xor (d271, d173, d179);
	nor (d272, d160, d174);
	nand (d273, d161, d176);
	nor (d274, d160, d163);
	and (d275, d177, d181);
	xnor (d276, d161, d169);
	xor (d277, d219, d269);
	or (d278, d231, d271);
	nor (d279, d242, d272);
	and (d280, d228, d260);
	or (d281, d242, d262);
	or (d282, d195, d245);
	xor (d283, d216, d264);
	nor (d284, d202, d267);
	nor (d285, d218);
	xnor (d286, d244, d259);
	xor (d287, d197, d246);
	buf (d288, d210);
	and (d289, d222, d272);
	buf (d290, d160);
	nor (d291, d190, d210);
	xnor (d292, d247, d264);
	xor (d293, d203, d241);
	or (d294, d219, d269);
	xor (d295, d206, d240);
	nand (d296, d210, d257);
	and (d297, d203, d270);
	xnor (d298, d256, d274);
	xnor (d299, d233, d273);
	xor (d300, d245, d271);
	nor (d301, d210, d249);
	buf (d302, d183);
	xor (d303, d211, d269);
	not (d304, d80);
	and (d305, d215);
	or (d306, d212, d274);
	xnor (d307, d191, d243);
	xor (d308, d246, d251);
	xor (d309, d206, d271);
	xnor (d310, d250, d257);
	and (d311, d199, d237);
	or (d312, d209, d267);
	not (d313, d141);
	not (d314, d213);
	xor (d315, d197, d248);
	or (d316, d188, d204);
	not (d317, d230);
	buf (d318, d190);
	xnor (d319, d201, d250);
	nor (d320, d209, d213);
	xor (d321, d208, d251);
	xor (d322, d189, d276);
	nor (d323, d195, d215);
	nand (d324, d202, d227);
	xnor (d325, d216, d259);
	xor (d326, d193, d197);
	nand (d327, d229, d272);
	and (d328, d190, d256);
	nand (d329, d264, d273);
	xor (d330, d236, d260);
	not (d331, d74);
	and (d332, d202, d267);
	xnor (d333, d202, d252);
	buf (d334, d239);
	not (d335, d151);
	nor (d336, d217, d225);
	xnor (d337, d250, d261);
	buf (d338, d146);
	buf (d339, d240);
	xor (d340, d210, d255);
	and (d341, d213, d215);
	or (d342, d201, d251);
	nor (d343, d233, d275);
	and (d344, d223, d249);
	buf (d345, d189);
	xnor (d346, d233, d257);
	buf (d347, d51);
	xor (d348, d215, d266);
	or (d349, d212, d243);
	or (d350, d205, d209);
	nand (d351, d207, d219);
	nor (d352, d203, d269);
	nor (d353, d225, d257);
	nand (d354, d216, d222);
	nand (d355, d228, d231);
	not (d356, d245);
	or (d357, d188, d255);
	xor (d358, d192, d195);
	nand (d359, d308, d324);
	nor (d360, d318, d345);
	xnor (d361, d348, d355);
	xnor (d362, d301, d323);
	or (d363, d315, d323);
	nand (d364, d288, d349);
	not (d365, d214);
	nand (d366, d300, d347);
	not (d367, d300);
	nand (d368, d312, d319);
	and (d369, d321, d333);
	xor (d370, d313, d334);
	or (d371, d283, d285);
	not (d372, d186);
	or (d373, d329, d337);
	or (d374, d297, d348);
	xor (d375, d324, d329);
	xnor (d376, d288, d293);
	not (d377, d192);
	nand (d378, d288, d328);
	or (d379, d342, d357);
	not (d380, d346);
	or (d381, d329, d356);
	buf (d382, d84);
	buf (d383, d354);
	xnor (d384, d295, d299);
	or (d385, d350, d354);
	and (d386, d313, d330);
	nand (d387, d328, d338);
	nor (d388, d292, d332);
	nor (d389, d332, d333);
	and (d390, d325, d351);
	or (d391, d279, d305);
	or (d392, d298, d340);
	or (d393, d283, d304);
	or (d394, d288, d355);
	buf (d395, d294);
	not (d396, d319);
	and (d397, d327, d357);
	xnor (d398, d291, d304);
	and (d399, d306, d313);
	nor (d400, d293, d310);
	xor (d401, d280, d289);
	assign f1 = d380;
	assign f2 = d397;
	assign f3 = d376;
	assign f4 = d365;
	assign f5 = d368;
	assign f6 = d387;
	assign f7 = d369;
	assign f8 = d376;
	assign f9 = d385;
	assign f10 = d375;
	assign f11 = d389;
	assign f12 = d359;
	assign f13 = d399;
	assign f14 = d387;
	assign f15 = d374;
	assign f16 = d367;
	assign f17 = d375;
	assign f18 = d372;
endmodule
