module CCGRCG5( x0, x1, f1, f2, f3, f4 );

	input x0, x1;
	output f1, f2, f3, f4;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252;

	buf (d1, x1);
	xor (d2, x1);
	and (d3, x0, x1);
	nor (d4, x1);
	xor (d5, x0);
	not (d6, x0);
	xnor (d7, x0, x1);
	xnor (d8, x0, x1);
	and (d9, x0, x1);
	xnor (d10, x1);
	nor (d11, x0, x1);
	xnor (d12, x0);
	nor (d13, x0);
	buf (d14, x0);
	xor (d15, x0, x1);
	nand (d16, x1);
	not (d17, x1);
	not (d18, d1);
	nor (d19, d9, d16);
	and (d20, d9, d16);
	nor (d21, d4, d11);
	not (d22, d6);
	xor (d23, d13, d17);
	and (d24, d10, d17);
	or (d25, d11, d12);
	xnor (d26, d1, d9);
	or (d27, d8, d17);
	or (d28, d2, d12);
	or (d29, d6, d7);
	xor (d30, d12, d13);
	buf (d31, d1);
	xnor (d32, d8, d15);
	nand (d33, d6, d14);
	xnor (d34, d3, d16);
	nand (d35, d3, d8);
	not (d36, d12);
	buf (d37, d9);
	buf (d38, d12);
	and (d39, d12, d15);
	nand (d40, d3, d5);
	nand (d41, d10, d15);
	nand (d42, d7, d14);
	xnor (d43, d9, d10);
	or (d44, d7, d13);
	xnor (d45, d4, d5);
	nand (d46, d2, d6);
	not (d47, d5);
	or (d48, d11);
	buf (d49, d4);
	xnor (d50, d2, d3);
	or (d51, d5, d10);
	buf (d52, d7);
	nand (d53, d2, d17);
	and (d54, d1, d2);
	xnor (d55, d3, d14);
	and (d56, d3, d15);
	and (d57, d7, d13);
	or (d58, d2, d8);
	or (d59, d4, d15);
	not (d60, d10);
	buf (d61, d11);
	xnor (d62, d7, d11);
	xnor (d63, d2, d13);
	nor (d64, d15);
	buf (d65, d17);
	and (d66, d12, d14);
	xor (d67, d7, d11);
	not (d68, d13);
	or (d69, d7, d12);
	xor (d70, d6, d12);
	or (d71, d1, d3);
	not (d72, d17);
	nand (d73, d2, d9);
	and (d74, d4, d8);
	nor (d75, d4, d12);
	buf (d76, d16);
	nor (d77, d2, d7);
	nand (d78, d1, d14);
	nor (d79, d15, d16);
	buf (d80, d6);
	or (d81, d1, d2);
	not (d82, d15);
	and (d83, d4, d13);
	nand (d84, d13, d16);
	or (d85, d68, d78);
	and (d86, d66, d81);
	and (d87, d27, d54);
	xnor (d88, d24, d45);
	buf (d89, d44);
	nand (d90, d31, d64);
	or (d91, d50, d60);
	nor (d92, d38, d43);
	or (d93, d61, d65);
	or (d94, d57, d60);
	buf (d95, d23);
	nand (d96, d60, d62);
	xnor (d97, d36, d50);
	or (d98, d62, d84);
	nand (d99, d79, d82);
	or (d100, d18, d30);
	xnor (d101, d54, d75);
	and (d102, d38, d49);
	xor (d103, d35, d76);
	nor (d104, d51, d55);
	nor (d105, d18, d54);
	xnor (d106, d45, d74);
	or (d107, d50, d53);
	nand (d108, d34, d68);
	buf (d109, d83);
	nor (d110, d28, d67);
	buf (d111, d14);
	nand (d112, d19, d24);
	xor (d113, d22, d46);
	and (d114, d58, d83);
	nand (d115, d48, d59);
	nor (d116, d58, d67);
	xor (d117, d47, d53);
	xnor (d118, d48, d53);
	buf (d119, d81);
	not (d120, d73);
	nand (d121, d41, d71);
	xnor (d122, d56, d73);
	and (d123, d26, d74);
	xnor (d124, d37, d80);
	xnor (d125, d56, d78);
	buf (d126, d52);
	not (d127, d84);
	xor (d128, d36, d67);
	and (d129, d41, d46);
	or (d130, d36, d44);
	nand (d131, d33, d35);
	xnor (d132, d36, d80);
	and (d133, d22, d61);
	or (d134, d38, d46);
	xor (d135, d57, d80);
	and (d136, d57, d78);
	or (d137, d49, d52);
	xor (d138, d36, d37);
	or (d139, d61, d74);
	not (d140, d49);
	xnor (d141, d46, d77);
	xnor (d142, d52, d77);
	xnor (d143, d25, d46);
	or (d144, d27, d35);
	xnor (d145, d23, d35);
	or (d146, d38, d71);
	or (d147, d53, d76);
	or (d148, d35, d67);
	xnor (d149, d28, d73);
	buf (d150, d64);
	xor (d151, d20, d79);
	buf (d152, d62);
	nor (d153, d37, d53);
	and (d154, d22, d69);
	nand (d155, d29, d32);
	xnor (d156, d52, d69);
	buf (d157, d54);
	xor (d158, d55, d67);
	xor (d159, d61, d74);
	xor (d160, d32, d53);
	not (d161, d66);
	xnor (d162, d146, d157);
	not (d163, d138);
	nand (d164, d106, d132);
	or (d165, d89, d142);
	nand (d166, d137, d145);
	buf (d167, d29);
	and (d168, d94, d108);
	xor (d169, d153, d154);
	nor (d170, d121, d147);
	xnor (d171, d99, d126);
	nor (d172, d122, d144);
	or (d173, d100, d121);
	xnor (d174, d128, d133);
	nand (d175, d98, d119);
	nor (d176, d91, d131);
	buf (d177, d61);
	and (d178, d117, d146);
	nor (d179, d98, d155);
	buf (d180, d49);
	or (d181, d92, d113);
	buf (d182, d136);
	not (d183, d9);
	or (d184, d110, d153);
	nor (d185, d105, d113);
	or (d186, d88, d98);
	xnor (d187, d92, d139);
	not (d188, d92);
	nor (d189, d85, d129);
	xor (d190, d124, d134);
	nor (d191, d88, d93);
	and (d192, d135, d153);
	xor (d193, d100, d114);
	or (d194, d87, d157);
	buf (d195, d100);
	and (d196, d96, d149);
	nand (d197, d115, d159);
	nor (d198, d110, d135);
	or (d199, d93, d121);
	buf (d200, d112);
	xor (d201, d113, d132);
	xor (d202, d109, d113);
	and (d203, d108, d127);
	xnor (d204, d132, d157);
	nor (d205, d98, d141);
	xor (d206, d124, d140);
	and (d207, d119, d144);
	nand (d208, d89);
	xnor (d209, d103, d110);
	buf (d210, d145);
	buf (d211, d86);
	and (d212, d141, d160);
	and (d213, d111, d117);
	nor (d214, d131, d147);
	nor (d215, d94, d135);
	xnor (d216, d85, d144);
	xor (d217, d97, d98);
	nand (d218, d131, d146);
	buf (d219, d124);
	nand (d220, d87, d93);
	nor (d221, d87, d119);
	or (d222, d105, d122);
	xor (d223, d86, d115);
	not (d224, d91);
	or (d225, d127, d152);
	or (d226, d141, d151);
	or (d227, d112, d136);
	not (d228, d56);
	xnor (d229, d89, d132);
	xor (d230, d104, d139);
	not (d231, d58);
	and (d232, d93, d100);
	not (d233, d125);
	xnor (d234, d129, d147);
	nand (d235, d90, d109);
	and (d236, d105, d147);
	or (d237, d110, d160);
	buf (d238, d111);
	xor (d239, d105, d117);
	and (d240, d106, d126);
	xnor (d241, d93, d96);
	or (d242, d97, d137);
	nor (d243, d106, d124);
	or (d244, d95, d138);
	nand (d245, d92, d133);
	xor (d246, d91, d128);
	xnor (d247, d120, d152);
	xor (d248, d135, d145);
	not (d249, d27);
	buf (d250, d38);
	nand (d251, d90, d123);
	not (d252, d135);
	assign f1 = d168;
	assign f2 = d177;
	assign f3 = d232;
	assign f4 = d162;
endmodule
