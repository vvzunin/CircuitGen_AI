module CCGRCG21( x0, x1, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12 );

	input x0, x1;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314, d315, d316, d317, d318, d319, d320, d321, d322, d323, d324, d325, d326, d327, d328, d329, d330, d331, d332, d333, d334, d335, d336, d337, d338, d339, d340, d341, d342, d343, d344, d345, d346, d347, d348, d349, d350, d351, d352, d353, d354, d355, d356, d357, d358, d359, d360, d361, d362, d363, d364, d365, d366, d367, d368, d369, d370, d371, d372, d373, d374, d375, d376, d377, d378, d379, d380, d381, d382, d383, d384, d385, d386, d387, d388, d389, d390, d391, d392, d393, d394, d395, d396, d397, d398, d399, d400, d401, d402, d403, d404, d405, d406, d407, d408, d409, d410, d411, d412, d413, d414, d415, d416, d417, d418, d419, d420, d421, d422, d423, d424, d425, d426, d427, d428;

	nand (d1, x0, x1);
	nor (d2, x1);
	nor (d3, x0);
	or (d4, x1);
	xor (d5, x0, x1);
	not (d6, x1);
	buf (d7, x1);
	nor (d8, x0, x1);
	nand (d9, x0, x1);
	xnor (d10, x0, x1);
	and (d11, x1);
	nand (d12, x0);
	xnor (d13, x0);
	and (d14, x0, x1);
	xnor (d15, x0, x1);
	buf (d16, x0);
	xor (d17, x0, x1);
	not (d18, x0);
	or (d19, x0);
	or (d20, x0, x1);
	xor (d21, x0);
	nor (d22, x0, x1);
	xor (d23, x1);
	and (d24, x0, x1);
	not (d25, d14);
	nor (d26, d1, d22);
	nand (d27, d9, d23);
	xor (d28, d6, d22);
	or (d29, d9, d14);
	or (d30, d2, d19);
	xor (d31, d15, d16);
	buf (d32, d11);
	buf (d33, d19);
	not (d34, d13);
	nand (d35, d1, d22);
	not (d36, d9);
	or (d37, d10, d20);
	and (d38, d9, d22);
	buf (d39, d17);
	nor (d40, d3, d14);
	nor (d41, d18, d24);
	xnor (d42, d2, d7);
	nor (d43, d7, d15);
	nand (d44, d1, d17);
	not (d45, d4);
	nor (d46, d7, d12);
	and (d47, d9, d24);
	buf (d48, d5);
	or (d49, d1, d3);
	xor (d50, d3, d5);
	buf (d51, d23);
	xnor (d52, d15, d23);
	or (d53, d9, d15);
	xnor (d54, d15, d16);
	or (d55, d1, d14);
	nand (d56, d1, d10);
	nor (d57, d2, d14);
	buf (d58, d3);
	or (d59, d23, d24);
	and (d60, d1, d11);
	and (d61, d2, d10);
	xnor (d62, d20, d24);
	not (d63, d24);
	xor (d64, d3, d12);
	and (d65, d7, d17);
	buf (d66, d7);
	and (d67, d21, d24);
	xnor (d68, d5, d10);
	xnor (d69, d23);
	xor (d70, d11, d18);
	buf (d71, d16);
	buf (d72, d12);
	xnor (d73, d5, d16);
	nor (d74, d1, d16);
	nand (d75, d6, d23);
	xnor (d76, d21, d23);
	and (d77, d6, d10);
	not (d78, d3);
	or (d79, d11, d16);
	and (d80, d1, d2);
	or (d81, d11, d22);
	xnor (d82, d1, d24);
	nor (d83, d6, d18);
	or (d84, d12, d13);
	xnor (d85, d10, d18);
	nand (d86, d2, d24);
	or (d87, d12, d18);
	buf (d88, d21);
	xnor (d89, d7, d22);
	xor (d90, d14, d17);
	nand (d91, d7, d11);
	and (d92, d7, d22);
	and (d93, d12, d15);
	xor (d94, d7, d14);
	xnor (d95, d10, d20);
	or (d96, d7, d14);
	buf (d97, d20);
	nand (d98, d35, d46);
	xor (d99, d30, d68);
	not (d100, d28);
	or (d101, d45, d80);
	xor (d102, d32, d62);
	not (d103, d1);
	nand (d104, d54, d65);
	and (d105, d60, d64);
	not (d106, d95);
	buf (d107, d89);
	or (d108, d66, d75);
	and (d109, d71, d78);
	xnor (d110, d76, d77);
	or (d111, d30, d57);
	not (d112, d74);
	nand (d113, d58, d67);
	nand (d114, d39, d47);
	not (d115, d72);
	xor (d116, d37, d69);
	or (d117, d57, d83);
	not (d118, d45);
	or (d119, d29, d75);
	xnor (d120, d73, d87);
	nor (d121, d65, d96);
	buf (d122, d77);
	or (d123, d76, d77);
	not (d124, d77);
	nand (d125, d34, d77);
	nand (d126, d52, d93);
	nor (d127, d53, d86);
	and (d128, d35, d80);
	nor (d129, d68, d78);
	buf (d130, d18);
	xnor (d131, d41, d77);
	nand (d132, d44, d54);
	buf (d133, d93);
	nand (d134, d77, d80);
	or (d135, d38, d88);
	xor (d136, d76);
	nor (d137, d48);
	not (d138, d80);
	and (d139, d31, d70);
	xor (d140, d75, d87);
	and (d141, d43, d75);
	and (d142, d55, d69);
	and (d143, d32, d49);
	xnor (d144, d67, d75);
	and (d145, d44, d80);
	nor (d146, d25, d92);
	xor (d147, d28, d96);
	not (d148, d94);
	buf (d149, d6);
	and (d150, d34, d89);
	xnor (d151, d40, d90);
	xnor (d152, d56, d68);
	xnor (d153, d32, d53);
	xor (d154, d92, d95);
	nor (d155, d25, d79);
	not (d156, d31);
	and (d157, d46, d57);
	nor (d158, d31);
	nand (d159, d70, d94);
	xor (d160, d25, d94);
	and (d161, d72, d89);
	and (d162, d51, d97);
	xor (d163, d60, d77);
	xor (d164, d43, d49);
	xnor (d165, d35, d36);
	xor (d166, d46, d93);
	xor (d167, d36, d68);
	nor (d168, d83, d95);
	buf (d169, d8);
	xnor (d170, d48, d73);
	nor (d171, d47, d48);
	nand (d172, d51, d68);
	xor (d173, d58, d66);
	buf (d174, d35);
	or (d175, d37, d97);
	and (d176, d65, d72);
	not (d177, d20);
	not (d178, d18);
	xnor (d179, d45, d75);
	xor (d180, d67, d68);
	buf (d181, d118);
	buf (d182, d156);
	nor (d183, d154, d179);
	xor (d184, d135, d155);
	not (d185, d104);
	xnor (d186, d142, d169);
	or (d187, d112);
	or (d188, d119, d152);
	nor (d189, d143, d150);
	or (d190, d105, d141);
	nand (d191, d105, d154);
	xor (d192, d100, d128);
	not (d193, d175);
	not (d194, d146);
	xnor (d195, d132, d147);
	buf (d196, d41);
	buf (d197, d160);
	nor (d198, d106, d172);
	and (d199, d142, d173);
	and (d200, d140, d164);
	nor (d201, d114, d134);
	or (d202, d119, d168);
	nor (d203, d102, d174);
	nor (d204, d128, d170);
	xor (d205, d116, d141);
	nand (d206, d121, d129);
	buf (d207, d92);
	buf (d208, d161);
	xnor (d209, d135, d161);
	not (d210, d65);
	xor (d211, d117, d132);
	or (d212, d123, d136);
	buf (d213, d121);
	or (d214, d118, d154);
	not (d215, d26);
	nand (d216, d100, d151);
	nor (d217, d109, d169);
	xor (d218, d112, d128);
	or (d219, d101, d131);
	buf (d220, d56);
	buf (d221, d204);
	buf (d222, d46);
	not (d223, d216);
	xnor (d224, d182, d219);
	xor (d225, d215, d217);
	xor (d226, d206, d215);
	or (d227, d202, d211);
	xnor (d228, d206, d212);
	not (d229, d190);
	nor (d230, d182, d195);
	not (d231, d122);
	nor (d232, d189, d206);
	xnor (d233, d200, d201);
	nor (d234, d184, d189);
	nor (d235, d201, d204);
	not (d236, d27);
	and (d237, d186, d191);
	nand (d238, d197, d207);
	nor (d239, d189, d194);
	nor (d240, d189, d199);
	buf (d241, d195);
	xor (d242, d186, d212);
	buf (d243, d150);
	xor (d244, d194, d208);
	or (d245, d183, d193);
	xor (d246, d187, d209);
	not (d247, d202);
	nand (d248, d193, d218);
	xnor (d249, d209);
	nand (d250, d195, d214);
	not (d251, d75);
	or (d252, d184, d185);
	and (d253, d191, d207);
	xnor (d254, d185, d205);
	or (d255, d226, d243);
	or (d256, d231, d241);
	xor (d257, d236, d254);
	xor (d258, d235, d251);
	not (d259, d51);
	and (d260, d225, d231);
	nor (d261, d225, d236);
	buf (d262, d246);
	or (d263, d225, d238);
	not (d264, d210);
	nor (d265, d246, d254);
	not (d266, d133);
	xnor (d267, d225, d239);
	or (d268, d228, d254);
	and (d269, d223, d249);
	and (d270, d221);
	xnor (d271, d237, d246);
	nand (d272, d230, d244);
	buf (d273, d67);
	xor (d274, d238, d246);
	xnor (d275, d225, d254);
	nor (d276, d221, d228);
	xnor (d277, d229, d236);
	and (d278, d244, d250);
	xnor (d279, d229, d233);
	and (d280, d243, d246);
	not (d281, d30);
	or (d282, d240, d246);
	buf (d283, d68);
	buf (d284, d29);
	and (d285, d223, d233);
	nor (d286, d225, d249);
	xor (d287, d221, d254);
	nor (d288, d238, d243);
	or (d289, d242, d243);
	or (d290, d220, d251);
	xor (d291, d222, d238);
	nand (d292, d233, d241);
	xnor (d293, d231, d249);
	nor (d294, d232, d238);
	not (d295, d149);
	and (d296, d228, d246);
	nor (d297, d230, d246);
	xor (d298, d220, d249);
	and (d299, d233, d254);
	buf (d300, d123);
	xor (d301, d220, d239);
	nand (d302, d220, d243);
	xnor (d303, d226, d243);
	nor (d304, d246, d250);
	or (d305, d245, d249);
	or (d306, d244, d246);
	nand (d307, d246, d253);
	and (d308, d224, d251);
	or (d309, d223, d224);
	not (d310, d162);
	or (d311, d233, d247);
	nor (d312, d222, d250);
	nor (d313, d223);
	not (d314, d252);
	xnor (d315, d225, d249);
	and (d316, d233, d250);
	buf (d317, d86);
	or (d318, d232, d252);
	and (d319, d224);
	nand (d320, d231, d236);
	not (d321, d206);
	nand (d322, d227, d230);
	and (d323, d226, d234);
	xor (d324, d242, d248);
	nor (d325, d223, d227);
	nor (d326, d226, d230);
	not (d327, d187);
	xor (d328, d235, d254);
	xnor (d329, d236, d249);
	xor (d330, d220, d248);
	nand (d331, d246, d250);
	nor (d332, d231, d232);
	nor (d333, d225, d226);
	nor (d334, d221, d241);
	buf (d335, d138);
	nand (d336, d278, d312);
	nand (d337, d274, d312);
	nor (d338, d258, d261);
	or (d339, d324, d331);
	buf (d340, d106);
	nand (d341, d300, d325);
	nand (d342, d297, d317);
	buf (d343, d292);
	buf (d344, d2);
	xnor (d345, d312, d327);
	and (d346, d318, d328);
	not (d347, d53);
	nor (d348, d258, d329);
	nor (d349, d261, d322);
	nand (d350, d289, d304);
	and (d351, d303, d318);
	xor (d352, d294, d333);
	buf (d353, d38);
	nand (d354, d316, d318);
	xnor (d355, d273, d292);
	and (d356, d293, d294);
	xor (d357, d296, d312);
	not (d358, d242);
	buf (d359, d215);
	buf (d360, d108);
	or (d361, d269, d327);
	xor (d362, d286);
	nand (d363, d300, d333);
	xnor (d364, d282, d319);
	and (d365, d288, d315);
	buf (d366, d314);
	nand (d367, d260, d286);
	or (d368, d262, d333);
	and (d369, d260, d297);
	nand (d370, d319, d333);
	not (d371, d304);
	not (d372, d276);
	xor (d373, d276, d304);
	nor (d374, d288, d319);
	not (d375, d110);
	xnor (d376, d281, d293);
	nand (d377, d255, d322);
	nor (d378, d274, d315);
	nand (d379, d280, d299);
	or (d380, d268, d323);
	and (d381, d303, d331);
	xnor (d382, d306);
	xnor (d383, d287, d324);
	buf (d384, d83);
	nor (d385, d285, d302);
	buf (d386, d54);
	xnor (d387, d279, d330);
	nand (d388, d255, d316);
	not (d389, d100);
	nor (d390, d293, d310);
	not (d391, d266);
	xor (d392, d295, d309);
	buf (d393, d174);
	xnor (d394, d298, d326);
	xnor (d395, d279, d303);
	nor (d396, d256, d311);
	xor (d397, d261, d321);
	xor (d398, d276, d335);
	xor (d399, d293, d318);
	and (d400, d274, d300);
	xor (d401, d273, d275);
	buf (d402, d228);
	not (d403, d253);
	and (d404, d303, d307);
	xnor (d405, d268, d272);
	not (d406, d200);
	nor (d407, d281, d322);
	and (d408, d260, d333);
	xor (d409, d281, d319);
	nor (d410, d318, d328);
	xor (d411, d284, d328);
	buf (d412, d142);
	xor (d413, d286, d292);
	nor (d414, d257, d264);
	xor (d415, d280, d289);
	nor (d416, d279, d324);
	nor (d417, d292, d310);
	nor (d418, d255, d294);
	buf (d419, d169);
	xor (d420, d257, d315);
	buf (d421, d304);
	nor (d422, d308, d328);
	and (d423, d264, d311);
	nor (d424, d258, d308);
	xnor (d425, d278, d318);
	xor (d426, d276, d279);
	xor (d427, d307, d320);
	nor (d428, d281, d315);
	assign f1 = d385;
	assign f2 = d407;
	assign f3 = d358;
	assign f4 = d382;
	assign f5 = d423;
	assign f6 = d403;
	assign f7 = d342;
	assign f8 = d410;
	assign f9 = d427;
	assign f10 = d342;
	assign f11 = d365;
	assign f12 = d407;
endmodule
