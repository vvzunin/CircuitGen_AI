module CCGRCG39( x0, x1, x2, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10 );

	input x0, x1, x2;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314;

	xor (d1, x1, x2);
	buf (d2, x2);
	or (d3, x0);
	xor (d4, x2);
	nand (d5, x2);
	buf (d6, x1);
	nand (d7, x0, x1);
	and (d8, x0, x1);
	and (d9, x1, x2);
	xor (d10, x0);
	nand (d11, x1, x2);
	and (d12, x0, x2);
	not (d13, x2);
	xnor (d14, x0, x1);
	or (d15, x1);
	nand (d16, x0, x2);
	buf (d17, x0);
	xor (d18, x0, x1);
	not (d19, x0);
	nand (d20, x1, x2);
	and (d21, x0, x1);
	and (d22, x0);
	or (d23, x0, x1);
	not (d24, x1);
	xor (d25, x0, x1);
	nand (d26, x0);
	nand (d27, x1);
	xnor (d28, x1);
	xnor (d29, x0, x2);
	nor (d30, x0, x1);
	xnor (d31, x1, x2);
	nor (d32, x0, x2);
	or (d33, x1, x2);
	or (d34, x0, x2);
	xnor (d35, x2);
	and (d36, x1, x2);
	and (d37, x2);
	and (d38, x0, x2);
	xnor (d39, x0, x2);
	nand (d40, x0, x1);
	nor (d41, x1, x2);
	xor (d42, x0, x2);
	nor (d43, x1);
	nor (d44, x2);
	xnor (d45, d15, d33);
	xor (d46, d23, d30);
	buf (d47, d23);
	xor (d48, d39, d42);
	buf (d49, d6);
	nand (d50, d4, d11);
	xor (d51, d24, d44);
	xnor (d52, d17, d38);
	and (d53, d22, d28);
	xor (d54, d2, d14);
	nand (d55, d30, d36);
	buf (d56, d30);
	or (d57, d27, d35);
	or (d58, d7, d17);
	not (d59, d33);
	or (d60, d15, d35);
	nor (d61, d6, d13);
	xnor (d62, d14, d26);
	nor (d63, d33, d36);
	and (d64, d4, d12);
	nand (d65, d9, d23);
	nor (d66, d14, d38);
	xor (d67, d27, d30);
	nor (d68, d17, d19);
	buf (d69, d21);
	buf (d70, d27);
	and (d71, d13, d20);
	not (d72, d7);
	nor (d73, d7, d12);
	nor (d74, d11, d22);
	not (d75, d20);
	nor (d76, d3, d25);
	and (d77, d18, d35);
	buf (d78, d4);
	xor (d79, d4, d7);
	buf (d80, d26);
	xor (d81, d33, d35);
	nand (d82, d7, d22);
	not (d83, d27);
	xor (d84, d2, d37);
	nand (d85, d40, d42);
	nor (d86, d3, d40);
	nor (d87, d19, d43);
	or (d88, d2, d23);
	buf (d89, d8);
	not (d90, d35);
	buf (d91, d43);
	not (d92, d28);
	or (d93, d9, d43);
	xor (d94, d6, d16);
	xnor (d95, d12, d26);
	nand (d96, d41, d43);
	and (d97, d3, d4);
	xnor (d98, d5, d37);
	not (d99, d32);
	nor (d100, d28, d35);
	not (d101, d13);
	nand (d102, d6, d25);
	nor (d103, d11, d30);
	or (d104, d15, d39);
	xor (d105, d6, d9);
	not (d106, d29);
	nor (d107, d14, d23);
	not (d108, d31);
	or (d109, d15, d34);
	xor (d110, d14, d15);
	nor (d111, d21, d30);
	buf (d112, d13);
	and (d113, d1, d30);
	or (d114, d18, d21);
	buf (d115, d36);
	and (d116, d9, d38);
	and (d117, d33, d41);
	or (d118, d9, d38);
	and (d119, d18, d27);
	buf (d120, d2);
	buf (d121, d18);
	and (d122, d25, d26);
	nand (d123, d29, d34);
	buf (d124, d9);
	buf (d125, d101);
	xor (d126, d53, d85);
	buf (d127, d65);
	and (d128, d75, d81);
	nand (d129, d70, d82);
	xor (d130, d48, d49);
	nand (d131, d85, d117);
	buf (d132, d74);
	and (d133, d57, d95);
	or (d134, d46, d99);
	nand (d135, d100, d101);
	xnor (d136, d80, d115);
	not (d137, d88);
	not (d138, d97);
	buf (d139, d108);
	nor (d140, d57, d121);
	buf (d141, d61);
	xnor (d142, d50, d78);
	xnor (d143, d83, d86);
	buf (d144, d49);
	nand (d145, d56, d59);
	or (d146, d47, d109);
	not (d147, d90);
	xnor (d148, d61, d78);
	not (d149, d52);
	buf (d150, d93);
	and (d151, d66);
	not (d152, d98);
	or (d153, d90, d101);
	not (d154, d108);
	or (d155, d118, d120);
	or (d156, d62, d75);
	and (d157, d68, d85);
	not (d158, d56);
	xor (d159, d46, d85);
	xnor (d160, d47, d99);
	xor (d161, d67, d107);
	or (d162, d88, d106);
	nand (d163, d85, d116);
	or (d164, d79, d101);
	xor (d165, d111, d114);
	or (d166, d66, d99);
	buf (d167, d54);
	xnor (d168, d65, d81);
	nand (d169, d51, d85);
	or (d170, d132, d143);
	buf (d171, d37);
	xor (d172, d143, d145);
	nor (d173, d133, d148);
	xnor (d174, d146, d152);
	nand (d175, d134, d154);
	not (d176, d16);
	and (d177, d151, d165);
	buf (d178, d69);
	and (d179, d136, d140);
	nand (d180, d137, d143);
	nor (d181, d140, d157);
	nand (d182, d127, d158);
	and (d183, d147, d150);
	or (d184, d152, d154);
	and (d185, d129, d140);
	nand (d186, d128, d153);
	nor (d187, d140, d166);
	buf (d188, d79);
	nor (d189, d138, d157);
	nor (d190, d156, d164);
	and (d191, d131, d143);
	not (d192, d59);
	and (d193, d140, d156);
	buf (d194, d83);
	xor (d195, d130, d160);
	xor (d196, d131, d164);
	buf (d197, d66);
	and (d198, d126, d162);
	xor (d199, d128, d131);
	buf (d200, d153);
	not (d201, d54);
	or (d202, d145, d162);
	xnor (d203, d129, d150);
	xnor (d204, d135, d142);
	buf (d205, d82);
	nand (d206, d142, d165);
	xnor (d207, d133, d134);
	and (d208, d131, d167);
	nand (d209, d157, d160);
	not (d210, d144);
	or (d211, d146, d166);
	nor (d212, d126, d155);
	and (d213, d134, d137);
	buf (d214, d156);
	xor (d215, d127, d134);
	buf (d216, d95);
	xnor (d217, d154, d160);
	nand (d218, d141, d156);
	or (d219, d130, d156);
	xor (d220, d160, d163);
	or (d221, d130, d152);
	and (d222, d132, d165);
	nor (d223, d146, d168);
	xor (d224, d129, d130);
	not (d225, d167);
	and (d226, d126, d160);
	nand (d227, d149, d166);
	xor (d228, d132, d141);
	or (d229, d134, d164);
	nand (d230, d130, d143);
	xnor (d231, d152, d168);
	not (d232, d101);
	nor (d233, d147, d148);
	or (d234, d144, d150);
	xnor (d235, d148, d159);
	xor (d236, d125, d161);
	not (d237, d232);
	xnor (d238, d173, d235);
	xor (d239, d201, d233);
	nor (d240, d172, d185);
	not (d241, d153);
	buf (d242, d128);
	buf (d243, d198);
	xnor (d244, d199, d206);
	nand (d245, d190, d209);
	nand (d246, d218, d220);
	xor (d247, d183, d189);
	xnor (d248, d228, d230);
	and (d249, d212, d213);
	xor (d250, d223, d233);
	nor (d251, d175, d190);
	nand (d252, d186, d222);
	buf (d253, d202);
	xnor (d254, d185, d216);
	or (d255, d174, d222);
	or (d256, d233, d236);
	or (d257, d192);
	xnor (d258, d171, d180);
	or (d259, d197, d223);
	not (d260, d15);
	nand (d261, d171, d187);
	not (d262, d93);
	nor (d263, d214, d225);
	or (d264, d173, d219);
	nor (d265, d202, d236);
	nor (d266, d197, d198);
	and (d267, d172, d195);
	nand (d268, d185, d220);
	not (d269, d163);
	nor (d270, d183, d232);
	and (d271, d206, d229);
	not (d272, d135);
	and (d273, d185, d188);
	xnor (d274, d175, d216);
	or (d275, d205, d228);
	buf (d276, d48);
	xor (d277, d179, d236);
	xnor (d278, d181, d182);
	or (d279, d208, d222);
	xor (d280, d195, d222);
	or (d281, d175, d229);
	nand (d282, d184, d215);
	not (d283, d61);
	buf (d284, d218);
	not (d285, d224);
	buf (d286, d131);
	nand (d287, d195, d199);
	nand (d288, d194, d218);
	and (d289, d179, d192);
	or (d290, d199, d235);
	nand (d291, d188, d221);
	or (d292, d176, d230);
	xor (d293, d175, d231);
	not (d294, d146);
	nand (d295, d174, d177);
	xor (d296, d187, d197);
	xnor (d297, d198, d232);
	or (d298, d205, d224);
	buf (d299, d199);
	and (d300, d181, d232);
	nor (d301, d174, d218);
	xor (d302, d191, d199);
	xnor (d303, d198, d219);
	or (d304, d173, d219);
	or (d305, d171, d207);
	or (d306, d178, d209);
	or (d307, d177, d213);
	xnor (d308, d196, d224);
	and (d309, d198, d224);
	nor (d310, d200, d222);
	nand (d311, d170, d211);
	nor (d312, d212, d233);
	xnor (d313, d200, d208);
	xnor (d314, d224, d234);
	assign f1 = d259;
	assign f2 = d262;
	assign f3 = d277;
	assign f4 = d255;
	assign f5 = d268;
	assign f6 = d242;
	assign f7 = d239;
	assign f8 = d288;
	assign f9 = d297;
	assign f10 = d286;
endmodule
