module CCGRCG115( x0, x1, x2, x3, x4, f1, f2 );

	input x0, x1, x2, x3, x4;
	output f1, f2;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314, d315, d316, d317, d318, d319, d320, d321, d322, d323, d324, d325, d326, d327, d328, d329, d330, d331, d332, d333, d334, d335, d336, d337, d338, d339, d340, d341, d342, d343, d344, d345, d346, d347, d348, d349, d350, d351, d352, d353, d354, d355, d356, d357, d358, d359, d360, d361, d362, d363, d364, d365, d366, d367, d368, d369, d370, d371, d372, d373, d374, d375, d376, d377, d378, d379, d380, d381, d382, d383, d384, d385, d386, d387, d388, d389, d390, d391, d392, d393, d394, d395, d396, d397, d398, d399;

	or (d1, x1, x4);
	buf (d2, x1);
	nor (d3, x1, x2);
	xor (d4, x2, x3);
	nor (d5, x0, x1);
	xnor (d6, x0, x2);
	xor (d7, x0, x1);
	or (d8, x0, x1);
	or (d9, x2);
	xor (d10, x1, x3);
	not (d11, x4);
	not (d12, x3);
	buf (d13, x0);
	nor (d14, x2, x4);
	not (d15, x1);
	xnor (d16, x0, x3);
	nor (d17, x4);
	nor (d18, d7, d10);
	and (d19, d4, d10);
	not (d20, d16);
	or (d21, d2, d10);
	and (d22, d6, d11);
	xnor (d23, d10, d13);
	nand (d24, d5);
	or (d25, d4, d14);
	not (d26, d11);
	xor (d27, d4, d5);
	not (d28, d15);
	nand (d29, d1, d9);
	xnor (d30, d5, d10);
	not (d31, d8);
	and (d32, d7, d11);
	xor (d33, d5, d12);
	and (d34, d1, d5);
	or (d35, d1);
	nor (d36, d9, d10);
	nand (d37, d4, d6);
	buf (d38, d13);
	xnor (d39, d9, d11);
	not (d40, d3);
	nor (d41, d2, d7);
	not (d42, d1);
	or (d43, d7, d17);
	nor (d44, d6, d14);
	xor (d45, d14, d15);
	or (d46, d8, d11);
	xnor (d47, d4, d8);
	and (d48, d4, d5);
	buf (d49, x3);
	not (d50, d12);
	nor (d51, d8, d11);
	not (d52, d9);
	nor (d53, d6, d10);
	buf (d54, x4);
	xor (d55, d8, d14);
	nand (d56, d1, d2);
	xor (d57, d6, d11);
	or (d58, d12);
	nor (d59, d8, d17);
	xnor (d60, d6, d17);
	xnor (d61, d3, d10);
	buf (d62, d11);
	nor (d63, d7, d11);
	nand (d64, d12, d17);
	or (d65, d5, d9);
	buf (d66, d4);
	or (d67, d3, d15);
	xor (d68, d31, d63);
	nand (d69, d21, d63);
	not (d70, d52);
	not (d71, d5);
	xor (d72, d41, d57);
	xor (d73, d25, d41);
	not (d74, d60);
	xor (d75, d53, d65);
	xor (d76, d30, d67);
	or (d77, d60);
	not (d78, d34);
	and (d79, d52, d59);
	not (d80, d6);
	and (d81, d53, d63);
	or (d82, d27, d58);
	not (d83, d2);
	not (d84, d36);
	buf (d85, d55);
	or (d86, d18, d54);
	not (d87, d66);
	xor (d88, d20, d57);
	buf (d89, d17);
	nor (d90, d20, d22);
	xnor (d91, d47, d51);
	buf (d92, d33);
	nand (d93, d32, d47);
	buf (d94, d63);
	nand (d95, d64, d67);
	not (d96, d26);
	buf (d97, d54);
	not (d98, d67);
	and (d99, d20, d58);
	buf (d100, d60);
	buf (d101, d31);
	nor (d102, d32, d61);
	xnor (d103, d24, d37);
	buf (d104, d29);
	nor (d105, d49, d55);
	nor (d106, d55, d63);
	not (d107, d37);
	nand (d108, d23, d57);
	not (d109, d55);
	nand (d110, d23, d67);
	xnor (d111, d34, d54);
	xnor (d112, d21, d22);
	nand (d113, d26, d56);
	buf (d114, d10);
	nand (d115, d24, d41);
	xnor (d116, d52, d66);
	xnor (d117, d27, d49);
	xnor (d118, d37, d58);
	and (d119, d23, d32);
	and (d120, d28, d36);
	and (d121, d23, d37);
	xnor (d122, d48, d60);
	xnor (d123, d24, d50);
	nor (d124, d27, d66);
	nand (d125, d37, d38);
	and (d126, d18, d34);
	and (d127, d29, d38);
	nor (d128, d18, d34);
	buf (d129, d34);
	xnor (d130, d33, d37);
	nor (d131, d20, d61);
	or (d132, d120, d129);
	and (d133, d68, d85);
	nand (d134, d98, d128);
	xnor (d135, d106, d127);
	xor (d136, d74, d75);
	nor (d137, d105, d126);
	xor (d138, d107, d120);
	xor (d139, d114, d120);
	buf (d140, d85);
	nor (d141, d81, d97);
	not (d142, d111);
	xor (d143, d87, d117);
	xor (d144, d93, d108);
	nand (d145, d79, d105);
	or (d146, d78, d81);
	nand (d147, d94, d103);
	nand (d148, d77, d129);
	nor (d149, d99, d110);
	xnor (d150, d69, d104);
	and (d151, d101, d115);
	or (d152, d96, d125);
	and (d153, d84, d123);
	xor (d154, d84, d104);
	buf (d155, d65);
	xnor (d156, d74, d129);
	xnor (d157, d75, d108);
	xor (d158, d70, d104);
	xor (d159, d89, d90);
	nand (d160, d93, d108);
	nand (d161, d79, d108);
	buf (d162, d71);
	buf (d163, d88);
	xor (d164, d89, d122);
	or (d165, d112);
	nor (d166, d114, d131);
	xor (d167, d99, d126);
	or (d168, d81, d110);
	xor (d169, d72, d99);
	nand (d170, d74, d100);
	xnor (d171, d137, d159);
	xnor (d172, d147, d167);
	nor (d173, d133, d154);
	nand (d174, d152, d159);
	buf (d175, d169);
	nand (d176, d155, d161);
	not (d177, d108);
	nand (d178, d155, d163);
	buf (d179, d87);
	nand (d180, d135, d152);
	not (d181, d119);
	nor (d182, d142, d152);
	and (d183, d141, d150);
	xor (d184, d143, d167);
	nand (d185, d135, d160);
	xnor (d186, d152, d164);
	nand (d187, d146, d152);
	and (d188, d133, d142);
	xnor (d189, d140, d152);
	xor (d190, d144, d166);
	nor (d191, d153, d168);
	xnor (d192, d150, d159);
	nor (d193, d152, d161);
	xor (d194, d144, d163);
	or (d195, d136, d141);
	xor (d196, d138, d169);
	or (d197, d140, d157);
	nor (d198, d151, d166);
	not (d199, d165);
	nor (d200, d157, d164);
	xor (d201, d151, d165);
	buf (d202, d74);
	buf (d203, d158);
	xnor (d204, d142, d160);
	buf (d205, d83);
	not (d206, d4);
	and (d207, d148, d168);
	or (d208, d136, d150);
	not (d209, d138);
	nand (d210, d138, d153);
	nand (d211, d135, d151);
	not (d212, d35);
	or (d213, d150, d156);
	xnor (d214, d133, d152);
	nand (d215, d144, d163);
	buf (d216, d96);
	xnor (d217, d142, d164);
	xnor (d218, d184, d189);
	and (d219, d187, d195);
	nand (d220, d175, d213);
	or (d221, d190, d208);
	and (d222, d187, d200);
	and (d223, d185, d194);
	not (d224, d123);
	nand (d225, d197, d204);
	nand (d226, d190, d206);
	xor (d227, d174, d192);
	xor (d228, d180, d185);
	and (d229, d187, d201);
	not (d230, d56);
	buf (d231, d135);
	xor (d232, d190, d195);
	or (d233, d195, d196);
	xnor (d234, d183, d186);
	xor (d235, d195, d208);
	and (d236, d194, d200);
	or (d237, d200, d207);
	xnor (d238, d198, d211);
	buf (d239, d152);
	xnor (d240, d213, d215);
	or (d241, d172, d199);
	xor (d242, d181, d193);
	and (d243, d184, d211);
	nand (d244, d181, d185);
	nand (d245, d172, d195);
	nand (d246, d203, d216);
	nand (d247, d177, d197);
	xnor (d248, d183, d184);
	nand (d249, d178, d179);
	xor (d250, d182, d183);
	xnor (d251, d200, d210);
	xor (d252, d192, d206);
	or (d253, d204, d216);
	xor (d254, d182, d198);
	xor (d255, d176, d206);
	xor (d256, d208, d217);
	xnor (d257, d197, d206);
	nor (d258, d177, d178);
	not (d259, d93);
	not (d260, d86);
	not (d261, d179);
	xor (d262, d174, d194);
	or (d263, d182, d199);
	xor (d264, d194, d195);
	xor (d265, d195, d196);
	xor (d266, d172, d182);
	nand (d267, d189, d210);
	and (d268, d180, d199);
	and (d269, d198, d204);
	xor (d270, d203, d211);
	xor (d271, d196, d206);
	not (d272, d200);
	and (d273, d174, d205);
	nand (d274, d201, d214);
	nor (d275, d178, d196);
	nor (d276, d190, d216);
	buf (d277, d86);
	or (d278, d177, d189);
	not (d279, d186);
	nor (d280, d171, d199);
	and (d281, d221, d267);
	and (d282, d237, d266);
	nor (d283, d226, d242);
	or (d284, d218, d249);
	and (d285, d265, d267);
	buf (d286, d111);
	buf (d287, d231);
	not (d288, d130);
	not (d289, d254);
	or (d290, d255, d269);
	nand (d291, d239, d254);
	xor (d292, d251, d268);
	xnor (d293, d221, d241);
	nand (d294, d236, d246);
	and (d295, d250, d267);
	xnor (d296, d261, d278);
	buf (d297, d143);
	buf (d298, d172);
	xor (d299, d234, d277);
	or (d300, d218, d243);
	or (d301, d227, d261);
	xnor (d302, d229, d265);
	xnor (d303, d240, d252);
	buf (d304, d27);
	not (d305, d256);
	xor (d306, d221, d231);
	xnor (d307, d236, d260);
	not (d308, d152);
	buf (d309, d175);
	or (d310, d251, d264);
	or (d311, d219, d266);
	buf (d312, d22);
	and (d313, d220, d230);
	not (d314, d155);
	nand (d315, d263);
	nor (d316, d235, d248);
	nand (d317, d230, d253);
	xnor (d318, d218, d278);
	not (d319, d229);
	or (d320, d261, d268);
	buf (d321, d247);
	buf (d322, d23);
	xor (d323, d244, d271);
	nand (d324, d246, d255);
	not (d325, d149);
	nor (d326, d236, d247);
	xnor (d327, d226, d269);
	xnor (d328, d230, d247);
	nand (d329, d228, d237);
	nor (d330, d235, d249);
	nand (d331, d233, d248);
	nor (d332, d219, d240);
	or (d333, d224, d258);
	and (d334, d243, d275);
	and (d335, d258, d273);
	nand (d336, d240);
	xnor (d337, d267, d270);
	not (d338, d31);
	and (d339, d227, d255);
	nor (d340, d224, d275);
	xnor (d341, d219, d229);
	buf (d342, d40);
	and (d343, d249, d271);
	xor (d344, d220, d235);
	nand (d345, d233, d258);
	nor (d346, d225, d247);
	xnor (d347, d221, d262);
	not (d348, d133);
	xnor (d349, d236, d238);
	or (d350, d220, d277);
	buf (d351, d72);
	nor (d352, d233, d247);
	nand (d353, d227, d257);
	nor (d354, d223, d266);
	nand (d355, d223, d252);
	buf (d356, d226);
	xor (d357, d222, d270);
	nor (d358, d224, d255);
	nor (d359, d254, d269);
	xnor (d360, d237, d259);
	or (d361, d253, d267);
	nor (d362, d255, d256);
	or (d363, d228, d258);
	nand (d364, d236, d260);
	or (d365, d219, d267);
	nand (d366, d284, d312);
	nand (d367, d286, d352);
	buf (d368, d20);
	nor (d369, d366);
	xor (d370, d366);
	not (d371, d281);
	nand (d372, d367, d368);
	buf (d373, d211);
	nor (d374, d368);
	buf (d375, d166);
	or (d376, d367);
	buf (d377, d326);
	not (d378, d65);
	or (d379, d366, d367);
	xor (d380, d366, d368);
	nand (d381, d367, d368);
	not (d382, d17);
	or (d383, d366, d367);
	nor (d384, d366, d368);
	or (d385, d366, d368);
	buf (d386, d296);
	not (d387, d310);
	not (d388, d89);
	not (d389, d296);
	nand (d390, d366, d368);
	not (d391, d105);
	and (d392, d366);
	nor (d393, d367, d368);
	nor (d394, d366, d368);
	and (d395, d367);
	and (d396, d367, d368);
	nand (d397, d366, d368);
	and (d398, d366, d368);
	xor (d399, d366, d367);
	assign f1 = d390;
	assign f2 = d399;
endmodule
