module CCGRCG142( x0, x1, x2, x3, x4, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16 );

	input x0, x1, x2, x3, x4;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314, d315, d316, d317, d318, d319, d320, d321, d322, d323, d324, d325, d326, d327, d328, d329, d330, d331, d332, d333, d334, d335, d336, d337, d338, d339, d340, d341, d342, d343, d344, d345, d346, d347, d348, d349, d350, d351, d352, d353, d354, d355, d356, d357, d358, d359, d360, d361, d362, d363, d364, d365, d366, d367, d368, d369, d370, d371, d372, d373, d374, d375, d376, d377, d378, d379, d380, d381, d382, d383, d384, d385, d386, d387, d388, d389, d390, d391, d392, d393, d394, d395, d396, d397, d398, d399, d400, d401, d402, d403;

	or (d1, x0, x2);
	and (d2, x1, x4);
	nand (d3, x3);
	xor (d4, x2, x3);
	xor (d5, x3, x4);
	xor (d6, x0);
	xor (d7, x1, x3);
	and (d8, x0, x3);
	and (d9, x1, x3);
	not (d10, x3);
	xnor (d11, x1, x3);
	xnor (d12, x1, x4);
	xor (d13, x0, x4);
	xnor (d14, x1);
	not (d15, x0);
	nor (d16, x0, x1);
	or (d17, x2, x3);
	or (d18, x4);
	or (d19, x3, x4);
	xor (d20, x2, x4);
	buf (d21, x4);
	buf (d22, x0);
	nand (d23, x2, x4);
	or (d24, x2, x3);
	xor (d25, x1, x2);
	not (d26, x2);
	and (d27, x2);
	and (d28, x0);
	or (d29, x0, x1);
	xnor (d30, x0, x1);
	nor (d31, x1, x3);
	or (d32, x1, x2);
	nor (d33, x0, x2);
	buf (d34, x3);
	and (d35, x0, x1);
	nand (d36, x1, x2);
	xor (d37, x1, x2);
	xnor (d38, x1, x2);
	xnor (d39, x1, x4);
	xnor (d40, x0, x2);
	nor (d41, x3, x4);
	buf (d42, x2);
	xor (d43, x3);
	xor (d44, x0, x2);
	or (d45, x3);
	not (d46, x4);
	nand (d47, x1, x4);
	or (d48, x2, x4);
	or (d49, d26, d29);
	xor (d50, d12, d41);
	or (d51, d38, d39);
	nor (d52, d31, d44);
	nor (d53, d15, d38);
	not (d54, d26);
	not (d55, d12);
	xor (d56, d4, d8);
	nand (d57, d2, d18);
	xnor (d58, d5, d47);
	or (d59, d23, d30);
	not (d60, d47);
	xnor (d61, d38, d47);
	not (d62, d50);
	nor (d63, d49, d52);
	and (d64, d55, d61);
	not (d65, d33);
	or (d66, d57, d58);
	and (d67, d52, d61);
	not (d68, d9);
	nor (d69, d50, d57);
	buf (d70, d46);
	nand (d71, d54, d55);
	not (d72, d17);
	buf (d73, d45);
	buf (d74, d20);
	xnor (d75, d49, d52);
	nor (d76, d55, d59);
	buf (d77, d52);
	xor (d78, d51, d54);
	xor (d79, d49, d61);
	and (d80, d61);
	or (d81, d51, d56);
	buf (d82, d25);
	xor (d83, d51, d56);
	nand (d84, d52, d59);
	nor (d85, d54, d57);
	buf (d86, d8);
	nor (d87, d52, d59);
	not (d88, d46);
	and (d89, d52, d53);
	xor (d90, d50, d58);
	xnor (d91, d50, d56);
	nand (d92, d53, d56);
	and (d93, d51, d59);
	buf (d94, d12);
	not (d95, d36);
	xor (d96, d55);
	buf (d97, d61);
	and (d98, d54, d61);
	nand (d99, d51, d52);
	or (d100, d54, d58);
	xor (d101, d49, d50);
	nand (d102, d52, d55);
	nor (d103, d62, d92);
	and (d104, d70, d73);
	not (d105, d78);
	not (d106, d68);
	and (d107, d64, d77);
	xnor (d108, d62, d82);
	nor (d109, d64, d93);
	not (d110, d63);
	xor (d111, d82, d92);
	not (d112, d34);
	xor (d113, d67, d83);
	nor (d114, d66, d81);
	nor (d115, d86, d91);
	and (d116, d89, d102);
	or (d117, d94, d100);
	buf (d118, d24);
	buf (d119, d60);
	nand (d120, d77, d81);
	buf (d121, d97);
	xnor (d122, d74, d91);
	buf (d123, d26);
	nor (d124, d88, d101);
	nand (d125, d67, d75);
	xor (d126, d94, d99);
	buf (d127, d64);
	and (d128, d77);
	nand (d129, d65, d68);
	and (d130, d64, d76);
	not (d131, d5);
	xnor (d132, d71, d79);
	not (d133, d98);
	xnor (d134, d79, d100);
	xor (d135, d97, d101);
	nand (d136, d68, d97);
	xnor (d137, d64, d88);
	nor (d138, d65, d90);
	xnor (d139, d72, d73);
	nor (d140, d71, d88);
	xor (d141, d81, d85);
	xnor (d142, d93, d95);
	and (d143, d66, d91);
	buf (d144, d18);
	nor (d145, d73, d78);
	xnor (d146, d85, d98);
	nand (d147, d92, d99);
	not (d148, d65);
	nand (d149, d70, d78);
	and (d150, d83, d94);
	and (d151, d70, d95);
	not (d152, d51);
	or (d153, d67, d90);
	xnor (d154, d64, d73);
	xor (d155, d72, d81);
	nand (d156, d68, d80);
	and (d157, d77, d93);
	nand (d158, d84, d87);
	or (d159, d86, d99);
	nor (d160, d98, d99);
	nor (d161, d66, d75);
	xnor (d162, d69, d86);
	nor (d163, d74, d84);
	xor (d164, d63, d79);
	nand (d165, d151, d159);
	nor (d166, d132, d139);
	buf (d167, d15);
	and (d168, d121, d138);
	nor (d169, d106, d146);
	xnor (d170, d122, d159);
	buf (d171, d94);
	not (d172, d123);
	nor (d173, d127, d153);
	xnor (d174, d122, d127);
	and (d175, d111, d140);
	nor (d176, d105, d142);
	buf (d177, d93);
	buf (d178, d145);
	nor (d179, d103, d155);
	nor (d180, d104, d133);
	buf (d181, d118);
	nor (d182, d135, d144);
	nand (d183, d131, d139);
	nor (d184, d156, d162);
	buf (d185, d17);
	nand (d186, d119, d134);
	buf (d187, d146);
	or (d188, d142);
	xnor (d189, d116, d122);
	xnor (d190, d111, d113);
	xor (d191, d131, d132);
	xor (d192, d124, d153);
	or (d193, d144, d145);
	nor (d194, d129, d162);
	xnor (d195, d105, d142);
	and (d196, d134, d149);
	nor (d197, d148, d162);
	or (d198, d111, d121);
	nor (d199, d120, d150);
	not (d200, d131);
	xnor (d201, d125, d160);
	or (d202, d107, d122);
	buf (d203, d73);
	xnor (d204, d155, d157);
	or (d205, d109, d163);
	or (d206, d116, d123);
	xor (d207, d103, d148);
	or (d208, d107, d145);
	buf (d209, d81);
	xnor (d210, d107, d153);
	xnor (d211, d111, d160);
	not (d212, d52);
	buf (d213, d154);
	or (d214, d125, d162);
	xnor (d215, d140, d142);
	and (d216, d138, d153);
	and (d217, d134, d137);
	or (d218, d134, d161);
	nand (d219, d113, d153);
	nand (d220, d122);
	nor (d221, d106, d134);
	xnor (d222, d106, d140);
	and (d223, d138, d147);
	xnor (d224, d139, d151);
	xnor (d225, d104, d120);
	nor (d226, d120, d132);
	xnor (d227, d138, d163);
	not (d228, d13);
	xnor (d229, d120, d134);
	or (d230, d139, d149);
	or (d231, d131, d162);
	nand (d232, d106, d164);
	nor (d233, d121, d143);
	nor (d234, d109, d136);
	or (d235, d109, d142);
	xor (d236, d107, d163);
	xnor (d237, d104, d155);
	xnor (d238, d109, d132);
	xor (d239, d109, d149);
	xnor (d240, d156, d162);
	xnor (d241, d131, d134);
	xnor (d242, d116, d153);
	nand (d243, d201, d214);
	xor (d244, d178, d236);
	not (d245, d15);
	xnor (d246, d165, d196);
	nor (d247, d187, d239);
	nand (d248, d193, d233);
	xnor (d249, d169, d191);
	nand (d250, d180, d182);
	nor (d251, d179, d199);
	and (d252, d196, d201);
	and (d253, d176, d214);
	xor (d254, d175, d217);
	nand (d255, d199, d237);
	nor (d256, d191, d215);
	nand (d257, d223, d240);
	not (d258, d188);
	not (d259, d148);
	or (d260, d176, d206);
	and (d261, d169, d240);
	and (d262, d167, d198);
	and (d263, d196, d214);
	or (d264, d201, d217);
	nand (d265, d194, d206);
	xor (d266, d174, d181);
	xor (d267, d169, d173);
	or (d268, d222, d234);
	buf (d269, d10);
	buf (d270, d109);
	not (d271, d259);
	nand (d272, d250, d259);
	nand (d273, d243, d253);
	nand (d274, d251, d255);
	buf (d275, d65);
	or (d276, d272, d273);
	and (d277, d272, d273);
	buf (d278, d112);
	and (d279, d271, d274);
	and (d280, d272, d274);
	xor (d281, d271);
	or (d282, d273, d274);
	and (d283, d272, d273);
	nor (d284, d271, d272);
	and (d285, d272);
	nor (d286, d271, d273);
	or (d287, d271, d272);
	and (d288, d273);
	xor (d289, d273, d274);
	buf (d290, d162);
	or (d291, d271, d273);
	buf (d292, d79);
	xor (d293, d271, d273);
	and (d294, d273, d274);
	and (d295, d272, d274);
	not (d296, d109);
	nor (d297, d272, d273);
	buf (d298, d75);
	and (d299, d271, d272);
	nor (d300, d274);
	not (d301, d116);
	and (d302, d271);
	or (d303, d273);
	or (d304, d272, d274);
	not (d305, d127);
	nor (d306, d271, d273);
	nand (d307, d273, d274);
	buf (d308, d11);
	not (d309, d48);
	not (d310, d223);
	xor (d311, d273, d274);
	or (d312, d272);
	buf (d313, d180);
	not (d314, d247);
	nor (d315, d304, d307);
	xnor (d316, d283, d295);
	or (d317, d290, d299);
	buf (d318, d156);
	nand (d319, d297, d299);
	and (d320, d301, d307);
	nor (d321, d279, d311);
	not (d322, d156);
	or (d323, d275, d295);
	xor (d324, d293, d300);
	xnor (d325, d297, d303);
	xor (d326, d296, d308);
	and (d327, d275, d284);
	nand (d328, d290, d305);
	or (d329, d284);
	or (d330, d285, d303);
	xnor (d331, d276, d309);
	not (d332, d174);
	nand (d333, d286, d300);
	xor (d334, d287, d290);
	xnor (d335, d294, d300);
	not (d336, d3);
	nand (d337, d299, d302);
	nor (d338, d285, d302);
	xnor (d339, d278, d287);
	xnor (d340, d288, d291);
	and (d341, d297, d299);
	and (d342, d279, d303);
	nor (d343, d305, d313);
	nand (d344, d292, d295);
	nor (d345, d285, d298);
	and (d346, d275, d300);
	xnor (d347, d293, d298);
	xor (d348, d281, d310);
	or (d349, d280, d306);
	buf (d350, d201);
	xor (d351, d285, d294);
	nand (d352, d278, d281);
	xor (d353, d287, d306);
	xnor (d354, d296, d304);
	not (d355, d133);
	and (d356, d278, d306);
	nand (d357, d276, d302);
	xnor (d358, d283, d289);
	and (d359, d283, d289);
	and (d360, d292, d295);
	not (d361, d280);
	xor (d362, d283, d302);
	or (d363, d296, d299);
	and (d364, d281, d300);
	xor (d365, d294, d309);
	buf (d366, d214);
	nor (d367, d280, d305);
	nor (d368, d305, d307);
	and (d369, d288, d290);
	xnor (d370, d291, d305);
	not (d371, d310);
	nor (d372, d335, d363);
	nand (d373, d341, d368);
	or (d374, d318, d344);
	nand (d375, d331, d369);
	not (d376, d264);
	xor (d377, d336, d338);
	or (d378, d320, d365);
	nand (d379, d316, d339);
	buf (d380, d318);
	nor (d381, d316, d332);
	not (d382, d178);
	nor (d383, d316, d328);
	or (d384, d314, d359);
	or (d385, d317, d364);
	xor (d386, d334, d362);
	not (d387, d243);
	nor (d388, d319, d333);
	nor (d389, d334, d367);
	xor (d390, d315, d352);
	xnor (d391, d316, d344);
	nand (d392, d322, d341);
	xnor (d393, d339, d370);
	or (d394, d342, d348);
	xnor (d395, d322, d334);
	buf (d396, d90);
	or (d397, d326, d345);
	buf (d398, d296);
	or (d399, d319, d364);
	xor (d400, d343);
	xor (d401, d337, d370);
	not (d402, d261);
	buf (d403, d106);
	assign f1 = d383;
	assign f2 = d387;
	assign f3 = d395;
	assign f4 = d375;
	assign f5 = d385;
	assign f6 = d403;
	assign f7 = d395;
	assign f8 = d403;
	assign f9 = d381;
	assign f10 = d384;
	assign f11 = d379;
	assign f12 = d372;
	assign f13 = d373;
	assign f14 = d391;
	assign f15 = d400;
	assign f16 = d390;
endmodule
