module CCGRCG149( x0, x1, x2, x3, x4, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17, f18, f19 );

	input x0, x1, x2, x3, x4;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17, f18, f19;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233;

	xnor (d1, x2, x4);
	not (d2, x1);
	and (d3, x2);
	nor (d4, x1, x3);
	or (d5, x0);
	and (d6, x0);
	xor (d7, x3);
	xor (d8, x1, x2);
	xor (d9, x2, x4);
	xor (d10, x0, x4);
	nand (d11, x0, x3);
	xnor (d12, x1);
	buf (d13, x2);
	xor (d14, x0, x1);
	xor (d15, x0);
	xnor (d16, x2);
	or (d17, x2, x3);
	xor (d18, x4);
	xor (d19, x0, x2);
	buf (d20, x4);
	nor (d21, x1, x4);
	nand (d22, x0, x4);
	nand (d23, x0, x1);
	nor (d24, x2);
	nand (d25, x4);
	buf (d26, x3);
	and (d27, x3, x4);
	and (d28, x1, x2);
	nand (d29, x1, x2);
	nand (d30, x3, x4);
	not (d31, x4);
	nand (d32, x0, x1);
	or (d33, x3, x4);
	xnor (d34, x0, x4);
	nand (d35, x0);
	buf (d36, x0);
	xnor (d37, x0, x1);
	or (d38, x1, x4);
	and (d39, x0, x4);
	xnor (d40, x3, x4);
	nand (d41, x0, x3);
	nor (d42, x0, x1);
	nor (d43, x0, x4);
	xnor (d44, x0, x1);
	xor (d45, x0, x1);
	and (d46, x3);
	or (d47, x0, x4);
	buf (d48, x1);
	not (d49, x0);
	nor (d50, x2, x4);
	nand (d51, x2, x3);
	nand (d52, x0, x2);
	and (d53, x0, x2);
	xor (d54, x1, x4);
	not (d55, x3);
	nor (d56, x1);
	nor (d57, x2, x3);
	nand (d58, x0, x2);
	xnor (d59, x1, x2);
	xnor (d60, x3, x4);
	nor (d61, x2, x4);
	xor (d62, x0, x4);
	xor (d63, x2, x3);
	or (d64, x0, x2);
	and (d65, x0, x2);
	xnor (d66, x2, x3);
	or (d67, d9, d11);
	or (d68, d15, d29);
	nand (d69, d15, d59);
	nand (d70, d25, d54);
	and (d71, d34, d40);
	or (d72, d42, d44);
	or (d73, d49, d57);
	xor (d74, d2, d10);
	buf (d75, d24);
	or (d76, d49, d64);
	xnor (d77, d11, d54);
	nand (d78, d17, d39);
	nand (d79, d4, d42);
	buf (d80, d64);
	xor (d81, d16, d65);
	buf (d82, d3);
	nor (d83, d22, d59);
	nor (d84, d37, d51);
	and (d85, d46, d61);
	not (d86, d53);
	xnor (d87, d13, d65);
	and (d88, d16, d24);
	nor (d89, d41, d49);
	or (d90, d8, d15);
	nand (d91, d26, d39);
	xor (d92, d48, d54);
	and (d93, d35, d59);
	xor (d94, d47, d58);
	or (d95, d21, d54);
	xnor (d96, d42, d62);
	and (d97, d33, d46);
	xor (d98, d16, d36);
	xnor (d99, d9, d38);
	or (d100, d36, d50);
	not (d101, d25);
	nand (d102, d9);
	or (d103, d9, d48);
	nor (d104, d16, d28);
	not (d105, d13);
	xor (d106, d30, d33);
	not (d107, d34);
	and (d108, d20, d40);
	and (d109, d42, d63);
	xor (d110, d17, d62);
	not (d111, d4);
	or (d112, d10, d36);
	not (d113, d61);
	xor (d114, d15, d35);
	or (d115, d47, d48);
	or (d116, d23, d27);
	xnor (d117, d50);
	and (d118, d25, d66);
	or (d119, d27, d36);
	nand (d120, d19, d53);
	nand (d121, d24, d26);
	xor (d122, d5, d66);
	nor (d123, d15, d21);
	not (d124, d35);
	xor (d125, d36, d60);
	xor (d126, d1, d52);
	not (d127, d28);
	and (d128, d4, d14);
	xnor (d129, d30, d36);
	nand (d130, d33, d49);
	or (d131, d7, d49);
	xnor (d132, d41, d63);
	nor (d133, d18, d55);
	xnor (d134, d14, d42);
	xnor (d135, d48, d60);
	xor (d136, d21, d28);
	nor (d137, d30, d51);
	nor (d138, d2, d39);
	xnor (d139, d3, d58);
	xnor (d140, d96, d117);
	xnor (d141, d74, d101);
	nand (d142, d72, d86);
	xor (d143, d111, d125);
	xor (d144, d70, d101);
	xor (d145, d90, d104);
	nand (d146, d86, d123);
	nand (d147, d68, d100);
	not (d148, d49);
	and (d149, d101, d106);
	xor (d150, d122, d128);
	buf (d151, d33);
	xnor (d152, d73, d134);
	nand (d153, d78, d91);
	buf (d154, d126);
	and (d155, d71, d98);
	xnor (d156, d75, d108);
	or (d157, d91, d118);
	xnor (d158, d83, d125);
	not (d159, d57);
	xor (d160, d105, d113);
	xnor (d161, d70, d121);
	xnor (d162, d87, d101);
	xnor (d163, d87, d104);
	xnor (d164, d88, d104);
	buf (d165, d57);
	and (d166, d100, d101);
	nor (d167, d114, d136);
	or (d168, d74, d120);
	nor (d169, d83, d137);
	nand (d170, d92, d129);
	nand (d171, d117, d132);
	nor (d172, d114, d119);
	or (d173, d121, d135);
	xnor (d174, d96, d131);
	nor (d175, d72, d87);
	nand (d176, d75, d97);
	nor (d177, d115, d116);
	buf (d178, d65);
	xor (d179, d101, d133);
	buf (d180, d92);
	xor (d181, d71, d85);
	xor (d182, d96, d130);
	xnor (d183, d114, d131);
	buf (d184, d37);
	nor (d185, d72, d73);
	xor (d186, d89, d128);
	nor (d187, d74, d113);
	xnor (d188, d105, d112);
	and (d189, d115, d118);
	or (d190, d89, d122);
	nor (d191, d79, d131);
	xnor (d192, d81, d112);
	buf (d193, d39);
	not (d194, d84);
	xor (d195, d98, d110);
	xnor (d196, d67, d112);
	xor (d197, d74, d121);
	and (d198, d87, d131);
	buf (d199, d71);
	and (d200, d85, d124);
	buf (d201, d32);
	and (d202, d80, d126);
	xor (d203, d78, d138);
	nor (d204, d73, d116);
	or (d205, d166, d179);
	xnor (d206, d194, d200);
	nor (d207, d166, d181);
	nor (d208, d166, d199);
	or (d209, d166, d202);
	nand (d210, d166, d190);
	nor (d211, d141, d180);
	not (d212, d203);
	nand (d213, d148, d182);
	buf (d214, d105);
	not (d215, d20);
	and (d216, d174, d183);
	not (d217, d204);
	xor (d218, d165, d172);
	and (d219, d177, d194);
	buf (d220, d139);
	nand (d221, d164, d204);
	xor (d222, d188, d204);
	not (d223, d5);
	nand (d224, d174, d181);
	xor (d225, d170, d176);
	or (d226, d182, d188);
	and (d227, d142, d190);
	and (d228, d143, d181);
	not (d229, d187);
	and (d230, d142, d155);
	and (d231, d160, d165);
	buf (d232, d168);
	and (d233, d188, d194);
	assign f1 = d220;
	assign f2 = d207;
	assign f3 = d207;
	assign f4 = d232;
	assign f5 = d220;
	assign f6 = d230;
	assign f7 = d233;
	assign f8 = d215;
	assign f9 = d212;
	assign f10 = d205;
	assign f11 = d221;
	assign f12 = d230;
	assign f13 = d221;
	assign f14 = d233;
	assign f15 = d229;
	assign f16 = d221;
	assign f17 = d213;
	assign f18 = d209;
	assign f19 = d219;
endmodule
