module CCGRCG48( x0, x1, x2, x3, f1, f2, f3, f4, f5 );

	input x0, x1, x2, x3;
	output f1, f2, f3, f4, f5;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99;

	buf (d1, x3);
	buf (d2, x0);
	not (d3, x2);
	or (d4, x2);
	xor (d5, x0, x1);
	not (d6, x0);
	nor (d7, x0, x3);
	nor (d8, x3);
	buf (d9, x2);
	xor (d10, x1);
	and (d11, x0, x1);
	buf (d12, x1);
	or (d13, x0, x1);
	xnor (d14, x2, x3);
	nand (d15, x2);
	nor (d16, x2, x3);
	xor (d17, x1, x2);
	xor (d18, x0, x1);
	and (d19, x1);
	and (d20, x0, x3);
	nand (d21, x2, x3);
	or (d22, x0, x2);
	not (d23, x3);
	nor (d24, x0, x2);
	and (d25, x1, x2);
	nor (d26, x1, x3);
	and (d27, x0, x2);
	nand (d28, x0, x1);
	xnor (d29, x2);
	or (d30, x0, x3);
	not (d31, x1);
	or (d32, x0, x3);
	nand (d33, x2, x3);
	nand (d34, x0);
	and (d35, x2, x3);
	not (d36, d8);
	buf (d37, d20);
	xnor (d38, d5, d35);
	xnor (d39, d5, d34);
	or (d40, d17, d20);
	not (d41, d5);
	and (d42, d5, d31);
	or (d43, d13);
	nand (d44, d19, d23);
	nor (d45, d11, d30);
	xnor (d46, d3, d7);
	buf (d47, d7);
	xor (d48, d18, d32);
	xor (d49, d4, d32);
	or (d50, d10, d29);
	or (d51, d25, d26);
	nor (d52, d10, d27);
	xor (d53, d13, d14);
	xor (d54, d15, d18);
	not (d55, d11);
	nor (d56, d5, d33);
	buf (d57, d35);
	not (d58, d35);
	xnor (d59, d14, d21);
	xnor (d60, d25, d26);
	nand (d61, d6, d24);
	buf (d62, d24);
	nor (d63, d53, d61);
	buf (d64, d59);
	and (d65, d38, d61);
	and (d66, d43, d61);
	buf (d67, d53);
	or (d68, d52, d55);
	nor (d69, d44, d45);
	and (d70, d43, d55);
	xnor (d71, d45, d47);
	or (d72, d37, d42);
	buf (d73, d38);
	xor (d74, d45, d61);
	xnor (d75, d45, d49);
	and (d76, d37, d60);
	nand (d77, d50, d61);
	xnor (d78, d51, d54);
	xnor (d79, d43, d52);
	buf (d80, d33);
	xor (d81, d40, d47);
	nor (d82, d41, d60);
	or (d83, d39, d58);
	not (d84, d12);
	nand (d85, d44, d61);
	xor (d86, d54, d55);
	or (d87, d48, d59);
	xnor (d88, d38, d58);
	xnor (d89, d43, d44);
	not (d90, d55);
	or (d91, d41, d60);
	or (d92, d61);
	and (d93, d42, d52);
	nand (d94, d44, d52);
	nor (d95, d50, d56);
	and (d96, d38, d56);
	xnor (d97, d57, d59);
	xor (d98, d50, d52);
	nand (d99, d43, d59);
	assign f1 = d83;
	assign f2 = d75;
	assign f3 = d86;
	assign f4 = d95;
	assign f5 = d79;
endmodule
