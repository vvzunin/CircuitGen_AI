module CCGRCG121( x0, x1, x2, x3, x4, f1, f2, f3, f4, f5 );

	input x0, x1, x2, x3, x4;
	output f1, f2, f3, f4, f5;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314, d315, d316, d317, d318, d319, d320, d321, d322, d323, d324, d325, d326, d327, d328, d329, d330, d331, d332, d333, d334, d335, d336, d337, d338, d339, d340, d341, d342, d343, d344, d345, d346, d347, d348, d349, d350, d351, d352, d353, d354, d355, d356, d357, d358, d359, d360, d361, d362, d363, d364, d365, d366, d367, d368, d369, d370, d371, d372, d373, d374, d375, d376, d377, d378, d379, d380, d381, d382, d383, d384, d385, d386, d387, d388, d389, d390, d391, d392, d393, d394, d395, d396, d397, d398, d399, d400, d401, d402, d403, d404, d405, d406, d407, d408, d409, d410, d411, d412, d413, d414, d415, d416, d417, d418, d419, d420, d421, d422, d423, d424, d425, d426, d427, d428, d429, d430, d431, d432, d433, d434, d435, d436, d437, d438, d439, d440, d441, d442, d443, d444, d445, d446, d447, d448, d449, d450, d451, d452, d453, d454, d455, d456, d457, d458, d459, d460, d461, d462, d463, d464, d465, d466, d467, d468, d469, d470, d471, d472, d473, d474, d475, d476, d477, d478, d479, d480, d481, d482, d483, d484, d485, d486, d487, d488, d489, d490, d491, d492, d493, d494, d495, d496;

	xor (d1, x1);
	xor (d2, x0, x4);
	not (d3, x3);
	buf (d4, x3);
	buf (d5, x1);
	xnor (d6, d2, d5);
	nand (d7, d3, d5);
	xor (d8, d2, d3);
	buf (d9, d1);
	and (d10, d6);
	nor (d11, d8);
	nor (d12, d6, d9);
	not (d13, x2);
	not (d14, d1);
	xor (d15, d7, d9);
	not (d16, d9);
	not (d17, d5);
	or (d18, d7, d9);
	xnor (d19, d8);
	xor (d20, d6, d8);
	not (d21, d6);
	nand (d22, d7);
	or (d23, d9);
	xor (d24, d6);
	xor (d25, d6, d9);
	nor (d26, d6, d7);
	nand (d27, d6, d9);
	or (d28, d6, d9);
	xor (d29, d8, d9);
	nor (d30, d6, d9);
	nand (d31, d8);
	or (d32, d6, d8);
	xnor (d33, d6, d9);
	not (d34, x0);
	xor (d35, d9);
	and (d36, d8, d9);
	or (d37, d6, d8);
	buf (d38, x4);
	xor (d39, d7, d8);
	nor (d40, d7, d8);
	xnor (d41, d6, d7);
	not (d42, d7);
	xor (d43, d8);
	not (d44, d3);
	xor (d45, d6, d8);
	not (d46, x1);
	xnor (d47, d6, d7);
	and (d48, d7, d9);
	nor (d49, d8, d9);
	nand (d50, d7, d9);
	nor (d51, d6, d8);
	and (d52, d6, d9);
	and (d53, d7, d8);
	and (d54, d6, d8);
	buf (d55, d7);
	or (d56, d20, d49);
	nor (d57, d23, d51);
	xor (d58, d36, d53);
	xnor (d59, d13, d20);
	and (d60, d37, d48);
	nor (d61, d41, d53);
	or (d62, d47, d49);
	or (d63, d31, d52);
	not (d64, d22);
	buf (d65, d22);
	nor (d66, d25, d33);
	and (d67, d24, d27);
	buf (d68, x2);
	nor (d69, d34, d49);
	nand (d70, d24, d41);
	xnor (d71, d52, d53);
	buf (d72, d49);
	not (d73, d11);
	xor (d74, d14, d47);
	not (d75, d47);
	and (d76, d22, d43);
	nand (d77, d26, d30);
	nand (d78, d30, d31);
	buf (d79, d48);
	nand (d80, d23, d24);
	not (d81, d44);
	xnor (d82, d33, d54);
	buf (d83, d46);
	not (d84, d25);
	or (d85, d26, d46);
	and (d86, d12, d52);
	or (d87, d35, d52);
	xor (d88, d13, d32);
	nor (d89, d33, d51);
	or (d90, d22, d45);
	nand (d91, d37, d42);
	nand (d92, d20, d28);
	nor (d93, d18, d44);
	buf (d94, d2);
	buf (d95, d32);
	buf (d96, d25);
	and (d97, d18, d38);
	nand (d98, d16, d31);
	buf (d99, x0);
	xor (d100, d10, d41);
	nand (d101, d16);
	nor (d102, d45, d47);
	not (d103, d15);
	not (d104, d52);
	and (d105, d44, d51);
	xnor (d106, d35, d51);
	xor (d107, d11, d20);
	xnor (d108, d34, d36);
	nand (d109, d12, d29);
	not (d110, d46);
	xor (d111, d40, d45);
	xnor (d112, d39, d52);
	xnor (d113, d19, d30);
	or (d114, d14, d29);
	buf (d115, d20);
	nor (d116, d24, d32);
	xnor (d117, d23, d37);
	not (d118, d18);
	nor (d119, d11, d42);
	nand (d120, d21, d42);
	or (d121, d18, d52);
	xor (d122, d13, d29);
	xnor (d123, d41);
	xor (d124, d13, d53);
	buf (d125, d50);
	xor (d126, d14, d49);
	xnor (d127, d10, d15);
	nor (d128, d10, d53);
	nand (d129, d27, d54);
	buf (d130, d42);
	or (d131, d17, d30);
	nand (d132, d10, d49);
	buf (d133, d4);
	not (d134, d105);
	and (d135, d66, d129);
	and (d136, d60, d77);
	xor (d137, d110, d118);
	xor (d138, d76, d106);
	nand (d139, d96, d121);
	not (d140, d31);
	xnor (d141, d104, d128);
	xnor (d142, d72, d106);
	xnor (d143, d84, d108);
	and (d144, d96, d117);
	nor (d145, d65, d74);
	nand (d146, d59, d71);
	xor (d147, d59, d70);
	buf (d148, d114);
	xor (d149, d78, d93);
	nand (d150, d69, d99);
	nand (d151, d87, d113);
	xor (d152, d77, d97);
	xor (d153, d98, d107);
	or (d154, d81, d130);
	not (d155, d29);
	and (d156, d74, d98);
	nor (d157, d103, d116);
	buf (d158, d5);
	xor (d159, d108, d120);
	and (d160, d58, d61);
	xor (d161, d88, d129);
	xnor (d162, d70);
	not (d163, d13);
	or (d164, d62);
	xnor (d165, d67, d131);
	and (d166, d81, d113);
	xnor (d167, d107, d126);
	xor (d168, d114, d120);
	nand (d169, d85, d96);
	nand (d170, d73, d113);
	xnor (d171, d56, d79);
	nand (d172, d71, d124);
	or (d173, d80, d113);
	nor (d174, d96, d103);
	not (d175, d62);
	nor (d176, d80, d124);
	buf (d177, d108);
	and (d178, d68, d93);
	or (d179, d64);
	not (d180, d118);
	xor (d181, d75, d117);
	nand (d182, d70, d128);
	buf (d183, d57);
	nand (d184, d60, d66);
	buf (d185, d76);
	not (d186, d42);
	nand (d187, d63, d84);
	not (d188, d32);
	nand (d189, d68, d84);
	xor (d190, d67, d119);
	nand (d191, d81, d86);
	xor (d192, d101, d120);
	xor (d193, d55, d69);
	nor (d194, d110, d122);
	buf (d195, d29);
	nand (d196, d117, d128);
	not (d197, d40);
	nand (d198, d81, d84);
	nand (d199, d81, d114);
	buf (d200, d111);
	and (d201, d72, d114);
	not (d202, d61);
	xnor (d203, d176, d193);
	xor (d204, d134, d150);
	and (d205, d140, d186);
	xnor (d206, d197, d201);
	xnor (d207, d139, d143);
	nand (d208, d149, d193);
	not (d209, d170);
	nor (d210, d156, d177);
	or (d211, d147, d194);
	or (d212, d163, d185);
	nand (d213, d149, d167);
	or (d214, d154, d180);
	xor (d215, d178, d193);
	not (d216, d163);
	xor (d217, d157, d201);
	xnor (d218, d140, d157);
	or (d219, d135, d165);
	or (d220, d160, d178);
	and (d221, d149, d153);
	nor (d222, d141, d191);
	xor (d223, d140, d153);
	and (d224, d151, d190);
	nand (d225, d136, d147);
	buf (d226, d193);
	nor (d227, d179, d199);
	or (d228, d144, d190);
	not (d229, d193);
	and (d230, d163, d201);
	buf (d231, d72);
	and (d232, d142, d146);
	xor (d233, d184, d185);
	and (d234, d145, d147);
	and (d235, d191, d193);
	not (d236, d161);
	not (d237, d50);
	nor (d238, d146, d168);
	or (d239, d173, d177);
	and (d240, d165, d181);
	xor (d241, d135, d186);
	buf (d242, d162);
	not (d243, d24);
	nand (d244, d190, d195);
	nor (d245, d152, d194);
	and (d246, d211, d220);
	or (d247, d209, d217);
	buf (d248, d129);
	buf (d249, d211);
	and (d250, d203, d238);
	nand (d251, d205, d213);
	xnor (d252, d236, d241);
	and (d253, d203, d223);
	nand (d254, d209, d215);
	xnor (d255, d207, d229);
	or (d256, d217, d244);
	buf (d257, d122);
	and (d258, d212, d223);
	or (d259, d202, d237);
	not (d260, d104);
	buf (d261, d149);
	nor (d262, d203, d207);
	nor (d263, d226, d237);
	nand (d264, d218, d226);
	buf (d265, d236);
	and (d266, d214, d235);
	not (d267, d156);
	xnor (d268, d224, d244);
	xor (d269, d230, d235);
	buf (d270, d243);
	buf (d271, d31);
	nor (d272, d206, d222);
	nand (d273, d202, d212);
	xor (d274, d207, d211);
	xnor (d275, d242, d243);
	or (d276, d241, d242);
	buf (d277, d96);
	not (d278, d88);
	not (d279, d214);
	xnor (d280, d205, d235);
	xor (d281, d206, d223);
	nor (d282, d202, d203);
	not (d283, d173);
	xnor (d284, d205, d241);
	buf (d285, d91);
	not (d286, d175);
	xor (d287, d206, d208);
	or (d288, d223, d245);
	nand (d289, d214, d225);
	xnor (d290, d211, d227);
	or (d291, d218, d237);
	not (d292, d79);
	and (d293, d234, d235);
	buf (d294, d13);
	xnor (d295, d207, d229);
	nand (d296, d217, d221);
	xor (d297, d228, d245);
	xor (d298, d214, d228);
	buf (d299, d205);
	xor (d300, d213, d241);
	not (d301, d160);
	not (d302, d201);
	nor (d303, d213, d214);
	xnor (d304, d212, d216);
	and (d305, d215, d225);
	or (d306, d206, d243);
	not (d307, d113);
	not (d308, d245);
	buf (d309, d242);
	xor (d310, d219, d227);
	or (d311, d202, d232);
	xor (d312, d221, d227);
	xnor (d313, d217, d241);
	not (d314, d34);
	nand (d315, d222, d229);
	buf (d316, d117);
	nand (d317, d267, d287);
	or (d318, d286, d311);
	or (d319, d260, d307);
	nor (d320, d296, d315);
	and (d321, d249, d296);
	or (d322, d300, d309);
	buf (d323, d165);
	xnor (d324, d257, d301);
	xnor (d325, d271, d277);
	xor (d326, d248, d255);
	or (d327, d251, d256);
	xor (d328, d250, d310);
	xnor (d329, d254, d292);
	xor (d330, d272, d276);
	not (d331, d314);
	xnor (d332, d285, d287);
	or (d333, d248, d261);
	not (d334, d194);
	or (d335, d253, d305);
	nor (d336, d294, d312);
	and (d337, d255, d292);
	nand (d338, d260, d262);
	xor (d339, d261, d310);
	nor (d340, d298, d302);
	nand (d341, d265, d316);
	xnor (d342, d287, d314);
	nand (d343, d319, d330);
	xor (d344, d336, d337);
	nor (d345, d322, d335);
	and (d346, d317, d322);
	xnor (d347, d320, d342);
	xor (d348, d318, d321);
	or (d349, d327, d338);
	or (d350, d322, d325);
	and (d351, d335, d340);
	xor (d352, d320, d327);
	nor (d353, d319, d333);
	not (d354, d184);
	xor (d355, d317, d341);
	nand (d356, d329, d334);
	and (d357, d318, d341);
	or (d358, d328, d334);
	nor (d359, d323, d325);
	or (d360, d323, d332);
	xnor (d361, d324, d335);
	xnor (d362, d321, d327);
	or (d363, d321, d329);
	or (d364, d326, d329);
	not (d365, d30);
	not (d366, d146);
	xor (d367, d322, d323);
	xor (d368, d320, d321);
	and (d369, d324, d338);
	xnor (d370, d327, d335);
	or (d371, d337, d342);
	and (d372, d328, d338);
	nand (d373, d322, d335);
	nand (d374, d319, d335);
	buf (d375, d75);
	nand (d376, d328, d342);
	not (d377, d155);
	xnor (d378, d318, d336);
	buf (d379, d63);
	nor (d380, d318, d326);
	buf (d381, d131);
	not (d382, d122);
	or (d383, d333);
	not (d384, d4);
	or (d385, d318, d325);
	and (d386, d325, d327);
	xnor (d387, d319, d337);
	and (d388, d328, d333);
	or (d389, d331, d340);
	xnor (d390, d333, d340);
	xor (d391, d324, d337);
	xnor (d392, d318, d326);
	xnor (d393, d320, d324);
	nor (d394, d320, d322);
	and (d395, d320, d321);
	nand (d396, d326, d331);
	xnor (d397, d325, d335);
	nand (d398, d338, d340);
	xor (d399, d320, d335);
	not (d400, d392);
	or (d401, d353, d362);
	or (d402, d380, d391);
	and (d403, d374, d389);
	not (d404, d140);
	xnor (d405, d348, d364);
	nand (d406, d363, d382);
	nor (d407, d347, d371);
	buf (d408, d369);
	nand (d409, d350, d389);
	nand (d410, d359, d362);
	xor (d411, d346, d350);
	nor (d412, d379, d396);
	or (d413, d393, d397);
	buf (d414, d386);
	xnor (d415, d346, d378);
	or (d416, d366, d384);
	and (d417, d358, d391);
	xnor (d418, d350, d369);
	and (d419, d345, d383);
	xor (d420, d353, d371);
	buf (d421, d343);
	nor (d422, d348, d349);
	not (d423, d281);
	not (d424, d190);
	xor (d425, d365, d383);
	xnor (d426, d354, d356);
	xnor (d427, d357, d399);
	nand (d428, d351, d376);
	nand (d429, d395, d397);
	buf (d430, d120);
	xor (d431, d369, d391);
	buf (d432, d278);
	not (d433, d251);
	xnor (d434, d361, d380);
	xor (d435, d383);
	or (d436, d346, d368);
	or (d437, d356, d392);
	and (d438, d347, d356);
	nand (d439, d366, d386);
	or (d440, d355, d384);
	nor (d441, d358, d391);
	xnor (d442, d369, d391);
	and (d443, d345, d366);
	not (d444, d394);
	nand (d445, d359, d380);
	nand (d446, d382, d393);
	nor (d447, d376, d377);
	not (d448, d103);
	nand (d449, d367, d389);
	not (d450, d296);
	xor (d451, d355, d360);
	xor (d452, d353, d398);
	and (d453, d358, d362);
	nor (d454, d344, d377);
	nor (d455, d375, d381);
	nor (d456, d380, d386);
	xor (d457, d386, d396);
	not (d458, d111);
	not (d459, d81);
	not (d460, d265);
	not (d461, d53);
	nor (d462, d375, d378);
	or (d463, d367, d388);
	or (d464, d380, d383);
	nand (d465, d347, d365);
	buf (d466, d143);
	xnor (d467, d391, d394);
	buf (d468, d389);
	nor (d469, d356, d398);
	xnor (d470, d386, d389);
	or (d471, d354, d379);
	buf (d472, d382);
	not (d473, d252);
	not (d474, d268);
	buf (d475, d146);
	xor (d476, d350, d383);
	nand (d477, d353, d357);
	xnor (d478, d378);
	and (d479, d345, d354);
	nand (d480, d375, d390);
	xor (d481, d385, d395);
	xor (d482, d349, d350);
	xnor (d483, d392, d399);
	or (d484, d369, d371);
	or (d485, d352, d374);
	not (d486, d12);
	or (d487, d368, d380);
	xor (d488, d357, d382);
	and (d489, d353, d356);
	nor (d490, d362, d398);
	not (d491, d322);
	not (d492, d35);
	not (d493, d206);
	buf (d494, d397);
	xor (d495, d355, d387);
	nand (d496, d353, d388);
	assign f1 = d495;
	assign f2 = d466;
	assign f3 = d436;
	assign f4 = d411;
	assign f5 = d436;
endmodule
