module CCGRCG31( x0, x1, x2, f1, f2, f3, f4, f5, f6 );

	input x0, x1, x2;
	output f1, f2, f3, f4, f5, f6;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143;

	nand (d1, x1, x2);
	buf (d2, x1);
	buf (d3, x2);
	xor (d4, x1, x2);
	not (d5, x0);
	or (d6, x0, x2);
	or (d7, x1);
	xor (d8, x0, x2);
	nand (d9, x2);
	not (d10, x1);
	and (d11, x1);
	nand (d12, x0, x2);
	or (d13, x0, x2);
	nand (d14, x1, x2);
	nor (d15, x0);
	and (d16, x0, x1);
	xor (d17, x1, x2);
	nor (d18, x0, x1);
	nand (d19, x0);
	xor (d20, x2);
	not (d21, x2);
	buf (d22, x0);
	or (d23, x0);
	and (d24, x0, x1);
	xor (d25, x0, x2);
	and (d26, x0);
	or (d27, x0, x1);
	and (d28, x1, x2);
	and (d29, x0, x2);
	or (d30, x2);
	xnor (d31, x0, x2);
	xnor (d32, x2);
	and (d33, x1, x2);
	xor (d34, x1);
	buf (d35, d32);
	nand (d36, d13, d22);
	buf (d37, d29);
	xor (d38, d9, d24);
	xor (d39, d4, d11);
	not (d40, d32);
	and (d41, d1, d3);
	xor (d42, d17, d19);
	buf (d43, d6);
	xor (d44, d8, d31);
	and (d45, d4, d24);
	xnor (d46, d9, d18);
	xor (d47, d8, d32);
	and (d48, d7, d26);
	xor (d49, d12, d22);
	not (d50, d10);
	nor (d51, d19, d31);
	xnor (d52, d29, d31);
	not (d53, d25);
	and (d54, d5, d7);
	nor (d55, d9, d19);
	xnor (d56, d8, d22);
	xnor (d57, d18, d33);
	xor (d58, d16, d19);
	or (d59, d8, d22);
	or (d60, d1, d24);
	buf (d61, d10);
	nor (d62, d16, d33);
	and (d63, d3, d17);
	nor (d64, d1, d8);
	and (d65, d4, d12);
	nor (d66, d14, d26);
	or (d67, d23, d25);
	and (d68, d13, d18);
	nand (d69, d18, d33);
	buf (d70, d9);
	not (d71, d18);
	or (d72, d8, d16);
	xnor (d73, d4, d23);
	xnor (d74, d12, d23);
	xor (d75, d5, d11);
	or (d76, d14);
	nor (d77, d12, d18);
	or (d78, d13, d17);
	xnor (d79, d21, d27);
	and (d80, d2, d12);
	or (d81, d27);
	and (d82, d20, d30);
	nor (d83, d1, d33);
	or (d84, d23, d34);
	xor (d85, d2, d7);
	buf (d86, d25);
	and (d87, d25, d28);
	xor (d88, d1, d4);
	xor (d89, d7, d15);
	xor (d90, d4, d21);
	and (d91, d1, d14);
	and (d92, d5, d10);
	and (d93, d19, d23);
	xnor (d94, d6, d24);
	nand (d95, d25, d26);
	xor (d96, d6, d24);
	and (d97, d3, d8);
	xor (d98, d15, d19);
	and (d99, d15, d22);
	nor (d100, d3, d27);
	xor (d101, d24, d28);
	buf (d102, d12);
	xor (d103, d4, d27);
	or (d104, d20, d33);
	xnor (d105, d6, d34);
	buf (d106, d15);
	nand (d107, d4, d13);
	or (d108, d6, d16);
	or (d109, d14, d26);
	buf (d110, d73);
	nor (d111, d41, d73);
	nand (d112, d110, d111);
	and (d113, d111);
	not (d114, d1);
	nor (d115, d111);
	nand (d116, d110);
	nor (d117, d110, d111);
	buf (d118, d108);
	xnor (d119, d110, d111);
	not (d120, d76);
	xor (d121, d110, d111);
	xor (d122, d110, d111);
	buf (d123, d69);
	xnor (d124, d110, d111);
	and (d125, d110, d111);
	nand (d126, d111);
	or (d127, d110, d111);
	nand (d128, d110, d111);
	nor (d129, d110);
	xnor (d130, d110);
	not (d131, d5);
	not (d132, d21);
	not (d133, d40);
	and (d134, d110, d111);
	buf (d135, d16);
	or (d136, d110);
	nor (d137, d110, d111);
	buf (d138, d30);
	buf (d139, d71);
	xor (d140, d110);
	xnor (d141, d111);
	not (d142, d55);
	not (d143, d4);
	assign f1 = d128;
	assign f2 = d142;
	assign f3 = d116;
	assign f4 = d113;
	assign f5 = d124;
	assign f6 = d123;
endmodule
