// Benchmark "CCGRCG74" written by ABC on Tue Feb 13 20:51:44 2024

module CCGRCG74 ( 
    x0, x1, x2,
    f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16,
    f17, f18, f19, f20  );
  input  x0, x1, x2;
  output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15,
    f16, f17, f18, f19, f20;
  wire new_n24_, new_n25_, new_n27_;
  assign new_n24_ = ~x0;
  assign new_n25_ = ~x1;
  assign f1 = ~x2 | ~new_n24_ | ~new_n25_;
  assign new_n27_ = ~x0 | ~x1;
  assign f2 = new_n27_ & (x0 | x2);
  assign f3 = ~new_n24_ | ~new_n25_;
  assign f4 = x2 & (x0 | x1);
  assign f5 = x2 & (x0 | x1);
  assign f6 = ~new_n24_ | ~new_n25_;
  assign f7 = x0;
  assign f8 = ~x2 | ~new_n24_ | ~new_n25_;
  assign f9 = x0;
  assign f10 = ~x2 | ~new_n24_ | ~new_n25_;
  assign f11 = ~x2 | ~new_n24_ | ~new_n25_;
  assign f12 = ~x2 | ~new_n24_ | ~new_n25_;
  assign f13 = x2 & (x0 | x1);
  assign f14 = ~x2 | ~new_n24_ | ~new_n25_;
  assign f15 = ~new_n24_ | ~new_n25_;
  assign f16 = x0;
  assign f17 = ~new_n24_ | ~new_n25_;
  assign f18 = new_n27_ & (x0 | x2);
  assign f19 = x0;
  assign f20 = ~x2 | ~new_n24_ | ~new_n25_;
endmodule


