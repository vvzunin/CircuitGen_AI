module CCGRCG65( x0, x1, x2, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15 );

	input x0, x1, x2;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157;

	and (d1, x0, x1);
	nand (d2, x2);
	nand (d3, x0, x1);
	nor (d4, x2);
	nand (d5, x0, x2);
	and (d6, x0);
	xor (d7, x0, x1);
	not (d8, x1);
	and (d9, x0, x1);
	xnor (d10, x0, x2);
	buf (d11, x1);
	xor (d12, x1, x2);
	xor (d13, x0, x2);
	or (d14, x1, x2);
	or (d15, x0, x1);
	and (d16, x0, x2);
	not (d17, x2);
	xnor (d18, x0);
	xnor (d19, x0, x1);
	xnor (d20, x1);
	xnor (d21, x2);
	buf (d22, x2);
	or (d23, x0);
	nand (d24, x0);
	nor (d25, x1, x2);
	not (d26, x0);
	and (d27, x2);
	nor (d28, x1);
	and (d29, x1);
	not (d30, d29);
	buf (d31, d26);
	or (d32, d4, d10);
	xor (d33, d6, d28);
	nand (d34, d1, d3);
	buf (d35, d4);
	or (d36, d3, d18);
	xor (d37, d4, d22);
	nand (d38, d3, d22);
	and (d39, d8, d17);
	buf (d40, d5);
	and (d41, d14, d29);
	nand (d42, d9, d22);
	and (d43, d2, d3);
	or (d44, d30, d40);
	nor (d45, d38, d42);
	nor (d46, d33, d35);
	xor (d47, d32, d34);
	nand (d48, d36, d40);
	nor (d49, d41, d42);
	buf (d50, d42);
	not (d51, d4);
	or (d52, d31, d36);
	nand (d53, d36, d42);
	buf (d54, d34);
	xor (d55, d36, d38);
	xor (d56, d37, d38);
	buf (d57, d11);
	xor (d58, d39, d43);
	buf (d59, d14);
	or (d60, d36, d37);
	xnor (d61, d37, d38);
	nand (d62, d31, d32);
	buf (d63, d30);
	xor (d64, d35, d37);
	or (d65, d33, d42);
	not (d66, d20);
	nor (d67, d34, d41);
	xor (d68, d33, d37);
	not (d69, d10);
	or (d70, d38, d43);
	buf (d71, d21);
	nand (d72, d31, d33);
	nand (d73, d39, d43);
	nor (d74, d35, d37);
	xor (d75, d31, d37);
	xor (d76, d30);
	not (d77, d35);
	xnor (d78, d52, d74);
	xnor (d79, d68, d76);
	or (d80, d47, d48);
	not (d81, d6);
	nand (d82, d68, d71);
	xor (d83, d56, d76);
	nand (d84, d55, d68);
	nor (d85, d65, d69);
	or (d86, d50, d59);
	and (d87, d64, d69);
	not (d88, d24);
	buf (d89, d54);
	xor (d90, d54, d63);
	or (d91, d62, d72);
	xor (d92, d61, d74);
	and (d93, d51, d54);
	not (d94, d11);
	not (d95, d63);
	or (d96, d63, d77);
	xnor (d97, d59, d77);
	or (d98, d48, d50);
	xor (d99, d57, d58);
	buf (d100, d40);
	nand (d101, d64, d68);
	or (d102, d52, d56);
	xnor (d103, d50, d53);
	and (d104, d58, d63);
	not (d105, d32);
	nand (d106, d70, d75);
	buf (d107, d29);
	nand (d108, d50, d63);
	nor (d109, d55, d65);
	buf (d110, d31);
	xor (d111, d56, d63);
	nor (d112, d47, d48);
	not (d113, d48);
	not (d114, d17);
	xor (d115, d64, d74);
	or (d116, d52, d59);
	not (d117, d74);
	not (d118, d50);
	and (d119, d57, d66);
	xnor (d120, d46, d76);
	nand (d121, d53, d62);
	buf (d122, d64);
	xor (d123, d54, d61);
	not (d124, d19);
	or (d125, d63, d71);
	xnor (d126, d61, d71);
	nor (d127, d47, d68);
	and (d128, d57, d68);
	nand (d129, d62, d72);
	and (d130, d46, d55);
	xnor (d131, d44, d51);
	buf (d132, x0);
	xor (d133, d66, d75);
	buf (d134, d19);
	nor (d135, d52, d55);
	xnor (d136, d54, d56);
	and (d137, d50, d77);
	xnor (d138, d49, d60);
	and (d139, d60, d73);
	xor (d140, d56, d57);
	and (d141, d59, d65);
	buf (d142, d55);
	nand (d143, d44, d59);
	nand (d144, d63, d74);
	xnor (d145, d62, d76);
	xor (d146, d52, d71);
	xor (d147, d50, d67);
	and (d148, d59, d74);
	nand (d149, d65, d66);
	and (d150, d45, d58);
	buf (d151, d76);
	and (d152, d75, d77);
	buf (d153, d27);
	nor (d154, d52, d57);
	buf (d155, d71);
	and (d156, d47, d62);
	xor (d157, d51, d75);
	assign f1 = d122;
	assign f2 = d92;
	assign f3 = d154;
	assign f4 = d156;
	assign f5 = d121;
	assign f6 = d102;
	assign f7 = d139;
	assign f8 = d126;
	assign f9 = d140;
	assign f10 = d151;
	assign f11 = d83;
	assign f12 = d134;
	assign f13 = d108;
	assign f14 = d116;
	assign f15 = d136;
endmodule
