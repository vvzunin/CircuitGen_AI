module CCGRCG71( x0, x1, x2, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17, f18 );

	input x0, x1, x2;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17, f18;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314, d315, d316, d317, d318, d319, d320, d321, d322, d323, d324, d325, d326, d327, d328, d329, d330, d331, d332, d333, d334, d335, d336, d337, d338, d339, d340, d341, d342, d343, d344, d345, d346, d347, d348, d349, d350, d351, d352, d353, d354, d355, d356, d357, d358, d359, d360, d361, d362, d363, d364, d365, d366, d367, d368, d369, d370, d371, d372, d373, d374, d375, d376, d377, d378, d379, d380, d381, d382, d383, d384, d385, d386, d387, d388, d389, d390, d391, d392, d393, d394, d395, d396, d397, d398, d399, d400, d401, d402, d403, d404, d405, d406, d407, d408, d409, d410, d411, d412, d413, d414, d415, d416, d417, d418, d419, d420, d421, d422, d423, d424, d425, d426, d427, d428, d429, d430, d431, d432, d433, d434, d435, d436, d437, d438, d439, d440, d441, d442, d443, d444, d445, d446, d447, d448, d449, d450, d451, d452, d453, d454, d455, d456, d457, d458, d459, d460, d461, d462, d463, d464, d465, d466, d467, d468, d469, d470, d471, d472, d473, d474, d475, d476, d477, d478, d479, d480, d481, d482, d483, d484, d485, d486, d487, d488, d489, d490, d491, d492, d493, d494, d495, d496, d497, d498, d499, d500, d501, d502, d503, d504, d505, d506, d507, d508, d509, d510, d511, d512, d513, d514, d515, d516, d517, d518, d519, d520, d521, d522, d523, d524, d525, d526, d527, d528, d529, d530, d531, d532, d533, d534, d535, d536, d537, d538, d539, d540, d541, d542, d543, d544, d545, d546, d547, d548, d549, d550;

	xor (d1, x0);
	or (d2, x0, x1);
	nand (d3, x0);
	nand (d4, x0, x2);
	xnor (d5, x0, x2);
	buf (d6, x1);
	buf (d7, x0);
	not (d8, x0);
	not (d9, x2);
	or (d10, x2);
	xor (d11, x1);
	nand (d12, x2);
	nor (d13, x0, x2);
	and (d14, x1, x2);
	xnor (d15, x0, x2);
	xor (d16, x2);
	nand (d17, x1, x2);
	not (d18, x1);
	or (d19, x0);
	nor (d20, x0, x2);
	xnor (d21, x0);
	nor (d22, x1);
	xor (d23, x0, x1);
	nor (d24, x0, x1);
	xor (d25, x0, x2);
	or (d26, x1, x2);
	and (d27, x0, x2);
	buf (d28, x2);
	xor (d29, x1, x2);
	nand (d30, x0, x2);
	or (d31, x1);
	xnor (d32, x1, x2);
	xnor (d33, x0, x1);
	nor (d34, x0);
	nor (d35, x0, x1);
	or (d36, d16, d30);
	xor (d37, d29, d34);
	not (d38, d11);
	buf (d39, d27);
	and (d40, d1, d5);
	nand (d41, d26);
	or (d42, d9, d26);
	xnor (d43, d13, d15);
	buf (d44, d28);
	xnor (d45, d1, d18);
	nand (d46, d17, d35);
	not (d47, d14);
	nor (d48, d14, d15);
	xor (d49, d12, d21);
	xnor (d50, d10, d16);
	and (d51, d5, d7);
	and (d52, d10, d29);
	and (d53, d28, d32);
	and (d54, d10, d21);
	nand (d55, d23, d30);
	xnor (d56, d12, d24);
	or (d57, d10, d31);
	and (d58, d15, d27);
	nor (d59, d20, d24);
	xnor (d60, d12, d21);
	and (d61, d8, d18);
	or (d62, d28, d30);
	nand (d63, d17, d24);
	nor (d64, d24, d29);
	and (d65, d2, d30);
	xnor (d66, d23, d35);
	not (d67, d2);
	not (d68, d9);
	nor (d69, d11, d22);
	nand (d70, d28, d33);
	nor (d71, d25, d35);
	xnor (d72, d7, d21);
	not (d73, d30);
	xnor (d74, d3, d13);
	nor (d75, d1, d12);
	nor (d76, d21, d35);
	xnor (d77, d10, d23);
	xor (d78, d6, d20);
	nor (d79, d15, d23);
	nor (d80, d2, d28);
	nor (d81, d14, d32);
	not (d82, d34);
	or (d83, d2, d32);
	xnor (d84, d2, d24);
	nor (d85, d20, d34);
	nand (d86, d18);
	or (d87, d9, d21);
	nand (d88, d22, d25);
	nor (d89, d5, d7);
	nand (d90, d27, d34);
	xor (d91, d16, d22);
	xnor (d92, d5, d20);
	xnor (d93, d8, d25);
	xnor (d94, d14, d22);
	nand (d95, d8, d21);
	nand (d96, d5, d15);
	xnor (d97, d23, d35);
	nand (d98, d26, d32);
	or (d99, d1, d26);
	buf (d100, d7);
	nor (d101, d7, d25);
	not (d102, d18);
	and (d103, d9, d22);
	or (d104, d16, d17);
	and (d105, d3, d21);
	nand (d106, d2, d29);
	nor (d107, d4, d32);
	and (d108, d13, d33);
	and (d109, d22, d24);
	not (d110, d26);
	and (d111, d33, d34);
	nand (d112, d4, d6);
	xor (d113, d5, d33);
	nand (d114, d4, d21);
	buf (d115, d3);
	nor (d116, d12, d25);
	buf (d117, d34);
	or (d118, d29, d31);
	nor (d119, d79, d112);
	nand (d120, d48, d98);
	buf (d121, d35);
	nand (d122, d76, d97);
	xnor (d123, d94, d103);
	nand (d124, d70, d86);
	xnor (d125, d40, d74);
	buf (d126, d85);
	nand (d127, d97, d104);
	and (d128, d43, d67);
	xnor (d129, d81, d115);
	or (d130, d83, d110);
	xnor (d131, d43, d114);
	or (d132, d71, d85);
	and (d133, d40, d58);
	buf (d134, d31);
	and (d135, d47, d79);
	not (d136, d70);
	buf (d137, d63);
	nor (d138, d44, d71);
	and (d139, d56, d60);
	or (d140, d89, d118);
	not (d141, d48);
	and (d142, d87, d107);
	not (d143, d59);
	not (d144, d92);
	buf (d145, d44);
	not (d146, d115);
	or (d147, d47, d107);
	nand (d148, d88);
	xor (d149, d72, d103);
	and (d150, d100, d106);
	buf (d151, d84);
	nor (d152, d40, d89);
	nand (d153, d82, d96);
	xor (d154, d47, d56);
	and (d155, d75, d91);
	xor (d156, d74, d81);
	nor (d157, d43, d63);
	xnor (d158, d74, d75);
	xor (d159, d64, d91);
	nand (d160, d108, d111);
	or (d161, d110, d116);
	buf (d162, d1);
	and (d163, d36, d97);
	xor (d164, d62, d108);
	not (d165, d77);
	nand (d166, d92, d112);
	xor (d167, d78, d98);
	buf (d168, d101);
	or (d169, d40, d77);
	buf (d170, d74);
	xor (d171, d86, d101);
	xnor (d172, d93, d101);
	buf (d173, d96);
	xnor (d174, d37, d118);
	nor (d175, d47, d108);
	buf (d176, d93);
	buf (d177, d51);
	buf (d178, d56);
	or (d179, d57, d92);
	xnor (d180, d59, d70);
	buf (d181, d8);
	buf (d182, d43);
	or (d183, d43, d49);
	nor (d184, d41, d95);
	xor (d185, d61, d110);
	xor (d186, d74, d89);
	nand (d187, d58, d77);
	or (d188, d41, d115);
	not (d189, d62);
	and (d190, d53, d117);
	nand (d191, d49, d105);
	or (d192, d58, d85);
	and (d193, d45, d67);
	buf (d194, d88);
	xnor (d195, d38, d84);
	buf (d196, d107);
	and (d197, d94, d110);
	buf (d198, d64);
	xnor (d199, d73, d100);
	or (d200, d36, d95);
	xor (d201, d93, d102);
	xnor (d202, d91, d97);
	not (d203, d78);
	nand (d204, d46, d52);
	and (d205, d57, d66);
	not (d206, d69);
	or (d207, d51, d90);
	xor (d208, d65, d79);
	xor (d209, d58, d100);
	or (d210, d92, d97);
	xnor (d211, d43, d116);
	or (d212, d145, d206);
	buf (d213, d135);
	xnor (d214, d121, d171);
	xnor (d215, d135, d142);
	or (d216, d126, d183);
	xnor (d217, d131, d191);
	and (d218, d145, d157);
	nand (d219, d180, d186);
	or (d220, d164, d194);
	and (d221, d142, d171);
	xor (d222, d170, d182);
	and (d223, d125, d200);
	xnor (d224, d163, d168);
	xor (d225, d145, d201);
	or (d226, d138, d139);
	not (d227, d199);
	xnor (d228, d121, d201);
	xnor (d229, d140, d203);
	or (d230, d120, d204);
	and (d231, d167, d207);
	and (d232, d164, d166);
	nor (d233, d123, d144);
	xnor (d234, d160, d173);
	xor (d235, d201, d207);
	nor (d236, d193, d197);
	nor (d237, d142, d191);
	not (d238, d134);
	buf (d239, d80);
	or (d240, d155, d158);
	nand (d241, d156, d202);
	or (d242, d166, d190);
	and (d243, d162, d167);
	xor (d244, d179, d194);
	nor (d245, d186, d195);
	or (d246, d227, d234);
	and (d247, d213, d237);
	or (d248, d220, d229);
	nor (d249, d219, d243);
	nor (d250, d237, d242);
	not (d251, d5);
	buf (d252, d123);
	xor (d253, d212, d215);
	and (d254, d212, d223);
	or (d255, d233, d244);
	buf (d256, d239);
	not (d257, d49);
	nor (d258, d213, d218);
	xor (d259, d220, d237);
	and (d260, d215, d222);
	xnor (d261, d223, d238);
	xnor (d262, d219, d220);
	xnor (d263, d232, d241);
	and (d264, d213, d214);
	nand (d265, d230, d235);
	or (d266, d230, d236);
	xnor (d267, d213, d244);
	xnor (d268, d224, d226);
	nor (d269, d222, d226);
	xor (d270, d230, d243);
	not (d271, d132);
	xnor (d272, d263, d265);
	buf (d273, d103);
	nand (d274, d249, d262);
	not (d275, d139);
	nor (d276, d262, d269);
	nor (d277, d256, d271);
	xnor (d278, d268, d269);
	nor (d279, d246, d266);
	nand (d280, d267, d269);
	or (d281, d255, d267);
	nand (d282, d246, d248);
	buf (d283, d175);
	nor (d284, d261, d268);
	xnor (d285, d249, d262);
	nor (d286, d261, d267);
	not (d287, d109);
	xnor (d288, d248, d266);
	or (d289, d265);
	not (d290, d80);
	nand (d291, d257, d271);
	nand (d292, d263, d271);
	nor (d293, d259);
	buf (d294, d258);
	xnor (d295, d260, d262);
	or (d296, d246, d269);
	xnor (d297, d256, d264);
	xnor (d298, d252, d262);
	xor (d299, d246, d265);
	xnor (d300, d251, d259);
	xnor (d301, d257, d258);
	buf (d302, d10);
	xor (d303, d256, d260);
	not (d304, d4);
	or (d305, d262, d267);
	nor (d306, d257, d269);
	xor (d307, d249, d250);
	xnor (d308, d258, d267);
	and (d309, d263, d267);
	or (d310, d246, d270);
	and (d311, d246, d254);
	buf (d312, d189);
	or (d313, d261);
	xor (d314, d256, d264);
	or (d315, d246, d258);
	nand (d316, d256, d265);
	buf (d317, d122);
	or (d318, d255, d269);
	buf (d319, d252);
	xor (d320, d248, d265);
	buf (d321, d222);
	nor (d322, d252, d269);
	buf (d323, d219);
	nor (d324, d252, d262);
	nor (d325, d253, d254);
	or (d326, d250, d261);
	xnor (d327, d256, d268);
	not (d328, d206);
	buf (d329, d128);
	buf (d330, d173);
	not (d331, d130);
	xor (d332, d255, d263);
	buf (d333, d95);
	nor (d334, d247, d257);
	xor (d335, d256, d271);
	nand (d336, d256, d257);
	nor (d337, d254, d260);
	xor (d338, d249, d268);
	buf (d339, d125);
	nor (d340, d246, d247);
	or (d341, d252, d256);
	nand (d342, d261, d262);
	or (d343, d252, d254);
	xnor (d344, d253, d268);
	not (d345, d50);
	nor (d346, d252, d261);
	xnor (d347, d262, d268);
	and (d348, d248, d267);
	and (d349, d259, d269);
	buf (d350, d259);
	and (d351, d257, d271);
	and (d352, d257, d266);
	buf (d353, d144);
	xnor (d354, d256, d271);
	and (d355, d248, d264);
	nor (d356, d246, d254);
	xnor (d357, d248, d254);
	buf (d358, d186);
	nand (d359, d265, d268);
	xor (d360, d250, d264);
	and (d361, d252, d271);
	xnor (d362, d248, d256);
	nor (d363, d251, d264);
	not (d364, d118);
	xor (d365, d247, d262);
	xnor (d366, d257, d270);
	nand (d367, d261, d271);
	nand (d368, d258, d269);
	buf (d369, d98);
	or (d370, d282, d285);
	not (d371, d274);
	buf (d372, d156);
	xnor (d373, d302, d339);
	not (d374, d47);
	buf (d375, d170);
	buf (d376, d369);
	xnor (d377, d285, d293);
	or (d378, d277, d345);
	and (d379, d300);
	not (d380, d299);
	nand (d381, d289, d341);
	buf (d382, d92);
	xor (d383, d293, d350);
	or (d384, d290, d362);
	nand (d385, d299, d307);
	and (d386, d373, d383);
	and (d387, d379, d382);
	nand (d388, d372, d383);
	buf (d389, d102);
	and (d390, d379, d384);
	nand (d391, d370, d379);
	xor (d392, d376, d383);
	nand (d393, d371, d375);
	nor (d394, d383, d384);
	not (d395, d236);
	nor (d396, d371, d377);
	not (d397, d200);
	xor (d398, d376, d377);
	buf (d399, d176);
	xnor (d400, d376, d378);
	nand (d401, d382, d384);
	not (d402, d12);
	nand (d403, d375, d379);
	nor (d404, d375, d380);
	or (d405, d376, d382);
	not (d406, d32);
	not (d407, d365);
	buf (d408, d70);
	xnor (d409, d382, d385);
	and (d410, d376, d380);
	and (d411, d373, d382);
	not (d412, d170);
	xor (d413, d383, d384);
	and (d414, d380, d383);
	and (d415, d371, d379);
	buf (d416, d19);
	nor (d417, d384, d385);
	nand (d418, d377, d381);
	and (d419, d371, d374);
	xor (d420, d375, d385);
	nor (d421, d372, d380);
	nand (d422, d371, d376);
	nand (d423, d380, d382);
	xor (d424, d372, d378);
	nor (d425, d403, d419);
	xnor (d426, d391, d420);
	not (d427, d347);
	xnor (d428, d390, d398);
	and (d429, d412, d417);
	not (d430, d352);
	nor (d431, d415, d418);
	buf (d432, d193);
	not (d433, d320);
	nor (d434, d417, d420);
	and (d435, d416, d419);
	or (d436, d396, d415);
	nor (d437, d386, d398);
	or (d438, d395, d423);
	or (d439, d395, d407);
	xor (d440, d393, d407);
	and (d441, d392, d420);
	nand (d442, d412, d420);
	not (d443, d172);
	xnor (d444, d406, d412);
	buf (d445, d330);
	buf (d446, d327);
	not (d447, d248);
	or (d448, d392, d401);
	nor (d449, d394, d422);
	or (d450, d396);
	or (d451, d402, d415);
	xnor (d452, d389, d409);
	xor (d453, d412, d424);
	nor (d454, d390);
	and (d455, d407, d408);
	and (d456, d403, d404);
	xor (d457, d410, d420);
	or (d458, d403, d422);
	or (d459, d389, d424);
	and (d460, d398, d404);
	buf (d461, d302);
	xnor (d462, d404);
	or (d463, d401, d408);
	nand (d464, d397, d410);
	nor (d465, d400, d412);
	or (d466, d393, d399);
	xnor (d467, d406, d420);
	xor (d468, d414, d424);
	or (d469, d404, d421);
	xnor (d470, d411, d418);
	not (d471, d213);
	not (d472, d98);
	xor (d473, d397, d408);
	and (d474, d386, d416);
	buf (d475, d223);
	nor (d476, d397, d409);
	xnor (d477, d389, d406);
	xnor (d478, d387, d421);
	nand (d479, d402, d407);
	xnor (d480, d398, d409);
	not (d481, d314);
	nand (d482, d401, d416);
	xor (d483, d407, d418);
	xnor (d484, d392, d407);
	not (d485, d343);
	nor (d486, d394, d421);
	not (d487, d111);
	nor (d488, d388, d396);
	and (d489, d399, d410);
	not (d490, d412);
	and (d491, d386, d399);
	and (d492, d410, d420);
	and (d493, d395, d411);
	xnor (d494, d387, d388);
	or (d495, d411, d413);
	or (d496, d386, d402);
	not (d497, d419);
	xnor (d498, d407, d424);
	or (d499, d404, d422);
	nand (d500, d399, d403);
	nand (d501, d392, d394);
	nor (d502, d453, d489);
	xor (d503, d455);
	buf (d504, d243);
	nor (d505, d449, d478);
	nor (d506, d444, d461);
	or (d507, d443, d479);
	nand (d508, d475, d480);
	not (d509, d387);
	or (d510, d439, d490);
	or (d511, d427, d449);
	not (d512, d104);
	nor (d513, d483, d497);
	or (d514, d442, d444);
	or (d515, d455, d491);
	not (d516, d384);
	not (d517, d329);
	xnor (d518, d438, d441);
	xor (d519, d439, d462);
	buf (d520, d108);
	buf (d521, d255);
	nand (d522, d430, d486);
	nor (d523, d435, d489);
	xnor (d524, d429, d489);
	xnor (d525, d436, d474);
	nand (d526, d445, d497);
	xnor (d527, d460, d475);
	xor (d528, d438, d461);
	nor (d529, d468, d470);
	nor (d530, d491, d498);
	and (d531, d442, d443);
	and (d532, d429, d494);
	xnor (d533, d465, d466);
	xnor (d534, d493, d501);
	not (d535, d8);
	nand (d536, d487, d494);
	xor (d537, d466, d480);
	xor (d538, d437, d478);
	xnor (d539, d466, d476);
	or (d540, d484, d496);
	xnor (d541, d433, d436);
	or (d542, d440, d454);
	not (d543, d351);
	nand (d544, d428, d501);
	and (d545, d438, d461);
	nor (d546, d476, d485);
	nor (d547, d428, d484);
	nand (d548, d452, d463);
	nand (d549, d488, d497);
	nand (d550, d431, d488);
	assign f1 = d514;
	assign f2 = d515;
	assign f3 = d536;
	assign f4 = d534;
	assign f5 = d548;
	assign f6 = d541;
	assign f7 = d523;
	assign f8 = d537;
	assign f9 = d537;
	assign f10 = d525;
	assign f11 = d540;
	assign f12 = d541;
	assign f13 = d510;
	assign f14 = d510;
	assign f15 = d513;
	assign f16 = d510;
	assign f17 = d542;
	assign f18 = d545;
endmodule
