module CCGRCG11( x0, x1, f1, f2, f3, f4, f5, f6, f7 );

	input x0, x1;
	output f1, f2, f3, f4, f5, f6, f7;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203;

	and (d1, x0, x1);
	or (d2, x0);
	nand (d3, x0, x1);
	xor (d4, x0, x1);
	buf (d5, x1);
	not (d6, x1);
	xnor (d7, x0);
	xor (d8, x0, x1);
	and (d9, x0, x1);
	xnor (d10, x0, x1);
	and (d11, x0);
	or (d12, x0, x1);
	buf (d13, x0);
	nand (d14, x0, x1);
	nand (d15, x0);
	not (d16, x0);
	and (d17, x1);
	or (d18, x1);
	xor (d19, x1);
	nand (d20, x1);
	nor (d21, x1);
	nor (d22, x0, x1);
	xnor (d23, x0, x1);
	nor (d24, x0, x1);
	xnor (d25, d13, d21);
	nor (d26, d4, d8);
	nor (d27, d13, d24);
	not (d28, d7);
	nand (d29, d2, d17);
	and (d30, d12, d13);
	xor (d31, d9, d17);
	nand (d32, d14, d22);
	buf (d33, d23);
	or (d34, d10, d17);
	not (d35, d23);
	xor (d36, d19, d20);
	or (d37, d12, d18);
	and (d38, d13, d16);
	nand (d39, d5, d14);
	not (d40, d8);
	xor (d41, d1, d3);
	nand (d42, d12, d22);
	and (d43, d14, d23);
	nor (d44, d22);
	nor (d45, d10, d16);
	not (d46, d21);
	nand (d47, d2, d13);
	xnor (d48, d5, d22);
	xor (d49, d12, d23);
	nand (d50, d3, d14);
	and (d51, d5, d11);
	xnor (d52, d10, d11);
	not (d53, d1);
	xnor (d54, d2, d20);
	buf (d55, d10);
	and (d56, d10, d18);
	xnor (d57, d7, d23);
	buf (d58, d6);
	xor (d59, d3, d19);
	and (d60, d7, d15);
	xnor (d61, d13, d20);
	xor (d62, d5, d13);
	xnor (d63, d3, d14);
	not (d64, d17);
	xor (d65, d2, d10);
	or (d66, d3, d10);
	xor (d67, d14, d24);
	xor (d68, d9, d22);
	xnor (d69, d3, d22);
	buf (d70, d3);
	not (d71, d22);
	nand (d72, d2, d3);
	or (d73, d14, d19);
	or (d74, d5, d17);
	and (d75, d13, d19);
	buf (d76, d8);
	or (d77, d11, d21);
	nand (d78, d5, d22);
	nand (d79, d2, d24);
	xnor (d80, d22, d23);
	or (d81, d20, d24);
	or (d82, d2, d3);
	xor (d83, d8, d16);
	and (d84, d1, d13);
	or (d85, d5, d17);
	xnor (d86, d14, d15);
	xnor (d87, d1, d12);
	nor (d88, d15, d16);
	xnor (d89, d8, d17);
	and (d90, d3, d4);
	nand (d91, d15, d18);
	or (d92, d10, d21);
	xor (d93, d13, d15);
	xor (d94, d15, d24);
	xnor (d95, d9, d15);
	nand (d96, d13, d19);
	xnor (d97, d11, d14);
	nand (d98, d3, d18);
	not (d99, d11);
	buf (d100, d20);
	xor (d101, d32, d54);
	nand (d102, d33, d77);
	xnor (d103, d44, d65);
	nor (d104, d58, d59);
	buf (d105, d74);
	xnor (d106, d51, d77);
	xor (d107, d74, d95);
	nor (d108, d75, d94);
	xnor (d109, d31, d73);
	xnor (d110, d34, d78);
	xnor (d111, d59, d97);
	xor (d112, d42, d56);
	nand (d113, d45, d91);
	and (d114, d36, d87);
	and (d115, d91);
	buf (d116, d1);
	not (d117, d35);
	not (d118, d27);
	not (d119, d20);
	buf (d120, d61);
	not (d121, d30);
	xnor (d122, d33, d88);
	nand (d123, d77, d91);
	or (d124, d30, d95);
	not (d125, d5);
	and (d126, d37, d99);
	xnor (d127, d49, d68);
	and (d128, d74, d90);
	nand (d129, d32, d70);
	xnor (d130, d32);
	not (d131, d12);
	xor (d132, d93, d94);
	nor (d133, d38, d89);
	not (d134, d25);
	not (d135, d38);
	xor (d136, d58, d89);
	buf (d137, d25);
	xor (d138, d44, d98);
	not (d139, d39);
	xor (d140, d47, d91);
	or (d141, d55, d66);
	and (d142, d37, d84);
	xnor (d143, d33, d52);
	or (d144, d78, d85);
	buf (d145, d64);
	nand (d146, d90);
	and (d147, d51, d58);
	and (d148, d58, d74);
	xor (d149, d37, d100);
	xnor (d150, d51, d99);
	or (d151, d48, d83);
	or (d152, d34, d77);
	or (d153, d26);
	buf (d154, d33);
	xor (d155, d73, d99);
	and (d156, d27, d65);
	xor (d157, d31, d66);
	xnor (d158, d73, d98);
	nand (d159, d27, d68);
	xor (d160, d58, d72);
	xnor (d161, d29, d34);
	nor (d162, d85);
	or (d163, d64, d94);
	or (d164, d42, d61);
	and (d165, d36, d99);
	xnor (d166, d57, d89);
	nand (d167, d42, d95);
	and (d168, d84, d88);
	xor (d169, d34, d42);
	or (d170, d46, d58);
	and (d171, d42, d90);
	and (d172, d95, d96);
	nand (d173, d51, d74);
	xor (d174, d64, d81);
	and (d175, d98, d99);
	not (d176, d72);
	not (d177, d55);
	not (d178, d50);
	or (d179, d36, d78);
	buf (d180, d97);
	and (d181, d54, d71);
	or (d182, d33, d58);
	and (d183, d61, d84);
	nor (d184, d62, d65);
	buf (d185, d183);
	nand (d186, d107, d108);
	and (d187, d185, d186);
	or (d188, d186);
	or (d189, d185);
	nand (d190, d185);
	buf (d191, d35);
	buf (d192, d48);
	and (d193, d185, d186);
	or (d194, d185, d186);
	xor (d195, d185, d186);
	nand (d196, d185, d186);
	nor (d197, d186);
	nand (d198, d186);
	buf (d199, d111);
	xor (d200, d186);
	nor (d201, d185, d186);
	xnor (d202, d185, d186);
	buf (d203, d155);
	assign f1 = d191;
	assign f2 = d192;
	assign f3 = d188;
	assign f4 = d190;
	assign f5 = d193;
	assign f6 = d198;
	assign f7 = d193;
endmodule
