module CCGRCG5( x0, x1, f1, f2, f3 );

	input x0, x1;
	output f1, f2, f3;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129;

	nor (d1, x0, x1);
	xnor (d2, x0, x1);
	nor (d3, x0, x1);
	or (d4, x1);
	xnor (d5, x0);
	buf (d6, x1);
	and (d7, x0, x1);
	nor (d8, x1);
	not (d9, x1);
	buf (d10, x0);
	xnor (d11, x1);
	nand (d12, x0, x1);
	not (d13, x0);
	xor (d14, x0, x1);
	and (d15, x0, x1);
	nand (d16, x0, x1);
	xnor (d17, x0, x1);
	and (d18, x1);
	or (d19, x0, x1);
	or (d20, x0, x1);
	xor (d21, x0, x1);
	nor (d22, x0);
	xor (d23, x1);
	nand (d24, x0);
	or (d25, x0);
	xor (d26, d11, d21);
	or (d27, d10, d21);
	nand (d28, d12, d19);
	nand (d29, d12, d17);
	buf (d30, d8);
	nor (d31, d2, d23);
	nand (d32, d8, d18);
	and (d33, d3, d19);
	xor (d34, d2, d19);
	xor (d35, d16, d22);
	xor (d36, d18, d22);
	not (d37, d13);
	buf (d38, d4);
	nand (d39, d4, d17);
	xor (d40, d32, d34);
	and (d41, d29, d38);
	buf (d42, d28);
	nand (d43, d27, d35);
	not (d44, d8);
	nor (d45, d26, d32);
	and (d46, d28, d37);
	xor (d47, d26, d38);
	buf (d48, d37);
	xor (d49, d30, d38);
	buf (d50, d33);
	buf (d51, d1);
	xnor (d52, d30, d38);
	xnor (d53, d26);
	and (d54, d46, d53);
	or (d55, d49, d53);
	not (d56, d12);
	xor (d57, d50, d51);
	xor (d58, d46, d48);
	nor (d59, d40, d45);
	nor (d60, d45);
	xnor (d61, d48, d50);
	and (d62, d41, d53);
	or (d63, d45, d49);
	not (d64, d35);
	and (d65, d40, d42);
	or (d66, d41, d52);
	not (d67, d50);
	xnor (d68, d40, d47);
	nand (d69, d44);
	xor (d70, d40, d53);
	or (d71, d45, d46);
	xnor (d72, d46, d52);
	nand (d73, d46, d52);
	or (d74, d44, d50);
	xor (d75, d42, d46);
	or (d76, d43, d52);
	nand (d77, d40, d47);
	nand (d78, d42, d49);
	and (d79, d45, d50);
	xnor (d80, d42, d48);
	xor (d81, d43, d48);
	buf (d82, d31);
	or (d83, d42, d50);
	and (d84, d44, d52);
	not (d85, d22);
	nor (d86, d48);
	nand (d87, d46, d48);
	xor (d88, d40, d42);
	not (d89, d24);
	nor (d90, d42, d49);
	xnor (d91, d42, d48);
	xnor (d92, d40, d50);
	nand (d93, d47, d52);
	and (d94, d41, d45);
	nand (d95, d40, d46);
	xor (d96, d41, d46);
	xnor (d97, d48, d49);
	xor (d98, d43, d45);
	or (d99, d42, d49);
	nor (d100, d48, d51);
	nor (d101, d43);
	nor (d102, d47, d48);
	nor (d103, d48, d51);
	xnor (d104, d40, d49);
	not (d105, d14);
	and (d106, d47, d48);
	xnor (d107, d41, d47);
	buf (d108, d46);
	xor (d109, d42, d47);
	xor (d110, d42);
	xnor (d111, d44, d49);
	and (d112, d46, d52);
	nor (d113, d40, d48);
	and (d114, d40, d41);
	xnor (d115, d46, d49);
	nor (d116, d40, d48);
	xor (d117, d43, d46);
	xnor (d118, d46, d47);
	xnor (d119, d43, d44);
	and (d120, d46, d47);
	and (d121, d48, d53);
	xnor (d122, d46, d49);
	or (d123, d43, d46);
	and (d124, d44, d50);
	xnor (d125, d42, d46);
	or (d126, d43, d50);
	or (d127, d50, d52);
	not (d128, d46);
	nor (d129, d45, d48);
	assign f1 = d65;
	assign f2 = d112;
	assign f3 = d98;
endmodule
