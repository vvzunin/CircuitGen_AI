module CCGRCG49( x0, x1, x2, x3, f1, f2, f3, f4, f5 );

	input x0, x1, x2, x3;
	output f1, f2, f3, f4, f5;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194;

	not (d1, x1);
	nand (d2, x0, x2);
	buf (d3, x2);
	nor (d4, x1, x2);
	xor (d5, x0, x1);
	or (d6, x1, x3);
	not (d7, x3);
	or (d8, x0, x1);
	xor (d9, x0, x1);
	xnor (d10, x2, x3);
	xnor (d11, x0, x2);
	buf (d12, x1);
	and (d13, x2, x3);
	xnor (d14, x1, x2);
	nand (d15, x0, x3);
	not (d16, x0);
	nand (d17, x1, x2);
	nor (d18, x1);
	nand (d19, x0);
	xnor (d20, x0, x1);
	and (d21, x0, x3);
	not (d22, x2);
	xor (d23, x1, x2);
	xnor (d24, x1);
	or (d25, x0, x3);
	nor (d26, x1, x3);
	and (d27, x1);
	nor (d28, x0, x1);
	or (d29, x2);
	nand (d30, x1, x3);
	and (d31, x2);
	or (d32, x1, x3);
	and (d33, x0, x2);
	xor (d34, x0, x3);
	buf (d35, x0);
	xor (d36, x0);
	nand (d37, x0, x2);
	or (d38, x1, x2);
	or (d39, x0, x3);
	nand (d40, x1);
	nor (d41, x3);
	and (d42, x0, x3);
	and (d43, x1, x2);
	nor (d44, x0);
	xor (d45, x0, x2);
	and (d46, x2, x3);
	xor (d47, x2, x3);
	nor (d48, x2);
	nor (d49, d11, d46);
	xnor (d50, d7, d47);
	buf (d51, d38);
	xnor (d52, d26, d32);
	nand (d53, d40, d46);
	buf (d54, d31);
	nor (d55, d13, d39);
	xor (d56, d32, d47);
	or (d57, d10, d48);
	nand (d58, d10, d29);
	and (d59, d10, d41);
	xor (d60, d32, d40);
	and (d61, d9, d26);
	not (d62, d33);
	nor (d63, d3, d45);
	and (d64, d16, d27);
	nand (d65, d2, d7);
	and (d66, d2, d13);
	nand (d67, d2, d34);
	xnor (d68, d18, d37);
	nor (d69, d35, d41);
	xor (d70, d43);
	nand (d71, d9, d42);
	nand (d72, d10, d32);
	nor (d73, d5, d46);
	buf (d74, d24);
	buf (d75, d32);
	not (d76, d24);
	and (d77, d3, d13);
	xor (d78, d21, d29);
	nand (d79, d36, d48);
	xor (d80, d31, d38);
	and (d81, d8, d41);
	xnor (d82, d37, d47);
	nand (d83, d25, d45);
	not (d84, d43);
	nand (d85, d44, d47);
	or (d86, d21, d45);
	or (d87, d16, d42);
	xnor (d88, d2, d34);
	xor (d89, d2, d27);
	xnor (d90, d6, d19);
	xnor (d91, d5, d19);
	xnor (d92, d6, d31);
	buf (d93, d4);
	buf (d94, d5);
	not (d95, d10);
	and (d96, d10, d47);
	xnor (d97, d28, d44);
	buf (d98, d13);
	or (d99, d27, d44);
	not (d100, d21);
	not (d101, d47);
	xnor (d102, d3, d30);
	not (d103, d30);
	xor (d104, d25, d30);
	not (d105, d1);
	nand (d106, d1, d42);
	xnor (d107, d32, d35);
	nor (d108, d33, d48);
	buf (d109, d17);
	or (d110, d14, d43);
	nand (d111, d8, d35);
	xor (d112, d13, d17);
	xor (d113, d19, d40);
	xor (d114, d1, d35);
	xnor (d115, d18, d38);
	nand (d116, d79, d88);
	nand (d117, d71, d99);
	buf (d118, d79);
	xnor (d119, d59, d103);
	or (d120, d51, d55);
	buf (d121, d92);
	xnor (d122, d72, d102);
	not (d123, d36);
	xor (d124, d102, d108);
	not (d125, d20);
	and (d126, d83, d100);
	nor (d127, d67, d79);
	not (d128, d72);
	xor (d129, d73, d97);
	nor (d130, d76, d85);
	xnor (d131, d70, d110);
	nor (d132, d67, d105);
	nand (d133, d100, d114);
	xor (d134, d64, d82);
	buf (d135, d33);
	and (d136, d81, d110);
	xnor (d137, d95, d97);
	buf (d138, d70);
	nor (d139, d71, d107);
	not (d140, d2);
	nor (d141, d122, d126);
	and (d142, d133, d138);
	or (d143, d127, d135);
	or (d144, d118, d127);
	buf (d145, d123);
	not (d146, d59);
	xor (d147, d134, d135);
	xor (d148, d122, d133);
	not (d149, d94);
	and (d150, d116, d126);
	not (d151, d98);
	or (d152, d119, d134);
	xor (d153, d121, d137);
	nor (d154, d135, d138);
	nand (d155, d125, d132);
	not (d156, d100);
	and (d157, d119, d121);
	not (d158, d138);
	nor (d159, d130, d132);
	and (d160, d118, d122);
	nand (d161, d121, d126);
	or (d162, d131, d134);
	nand (d163, d122, d134);
	xor (d164, d119, d121);
	and (d165, d122, d134);
	and (d166, d127, d135);
	nand (d167, d127, d137);
	nand (d168, d130, d131);
	xor (d169, d121, d126);
	xor (d170, d122, d126);
	xor (d171, d123, d125);
	or (d172, d116, d120);
	nor (d173, d120, d134);
	not (d174, d66);
	xor (d175, d118, d119);
	nand (d176, d125, d128);
	buf (d177, d2);
	xor (d178, d120, d130);
	xor (d179, d122, d138);
	or (d180, d118, d132);
	nor (d181, d124, d133);
	xor (d182, d117, d132);
	xnor (d183, d130, d131);
	xor (d184, d123, d126);
	not (d185, d89);
	buf (d186, d62);
	xnor (d187, d129, d136);
	xnor (d188, d120, d125);
	buf (d189, d78);
	nand (d190, d116, d127);
	nand (d191, d118, d125);
	xor (d192, d116, d139);
	nand (d193, d121, d123);
	xnor (d194, d120, d130);
	assign f1 = d186;
	assign f2 = d190;
	assign f3 = d156;
	assign f4 = d193;
	assign f5 = d183;
endmodule
