module CCGRCG55( x0, x1, x2, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10 );

	input x0, x1, x2;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299;

	nand (d1, x0, x2);
	or (d2, x1);
	nand (d3, x0, x1);
	and (d4, x1);
	nand (d5, x0, x2);
	not (d6, x1);
	and (d7, x1, x2);
	buf (d8, x0);
	nand (d9, x1);
	xnor (d10, x1);
	nor (d11, x1);
	or (d12, d9, d10);
	or (d13, d4, d11);
	or (d14, d3, d11);
	buf (d15, d4);
	or (d16, d3, d10);
	nand (d17, d1, d5);
	nand (d18, d1, d4);
	xnor (d19, d2, d4);
	or (d20, d6, d11);
	nand (d21, d10, d11);
	not (d22, x2);
	not (d23, d2);
	xnor (d24, d1, d8);
	not (d25, x0);
	xor (d26, d5);
	xnor (d27, d3, d11);
	nand (d28, d3, d7);
	not (d29, d1);
	and (d30, d3, d5);
	xnor (d31, d3, d9);
	and (d32, d6, d10);
	nor (d33, d7);
	nor (d34, d10, d11);
	and (d35, d2, d9);
	xnor (d36, d1, d7);
	xor (d37, d4);
	nand (d38, d2, d5);
	not (d39, d10);
	or (d40, d4);
	xnor (d41, d3, d10);
	nor (d42, d5, d7);
	not (d43, d8);
	buf (d44, d2);
	and (d45, d8, d11);
	and (d46, d3, d4);
	nor (d47, d3, d9);
	and (d48, d7);
	nor (d49, d2, d7);
	nand (d50, d5, d7);
	and (d51, d8, d9);
	nor (d52, d5, d10);
	and (d53, d7, d8);
	nor (d54, d2, d11);
	nand (d55, d6, d7);
	nand (d56, d4, d5);
	nor (d57, d2, d11);
	buf (d58, x2);
	buf (d59, d1);
	and (d60, d1, d9);
	nand (d61, d6);
	xor (d62, d8, d10);
	buf (d63, d7);
	xnor (d64, d6, d11);
	xor (d65, d2, d9);
	buf (d66, d6);
	xor (d67, d3, d7);
	and (d68, d3, d9);
	not (d69, d4);
	and (d70, d4, d6);
	nand (d71, d28, d70);
	xnor (d72, d29, d54);
	and (d73, d31, d65);
	nor (d74, d48, d54);
	and (d75, d16, d39);
	or (d76, d34, d50);
	nor (d77, d38, d49);
	not (d78, d18);
	or (d79, d21, d56);
	and (d80, d50, d57);
	xor (d81, d33, d45);
	not (d82, d68);
	nor (d83, d32, d38);
	or (d84, d44, d69);
	buf (d85, d16);
	xor (d86, d23, d56);
	xor (d87, d28, d36);
	nor (d88, d26, d66);
	not (d89, d58);
	xnor (d90, d14, d53);
	nor (d91, d60, d67);
	or (d92, d37, d41);
	xnor (d93, d37, d42);
	xor (d94, d14, d68);
	nor (d95, d65, d69);
	xnor (d96, d56, d68);
	nand (d97, d46, d57);
	and (d98, d19, d37);
	xor (d99, d14, d44);
	nor (d100, d28, d68);
	and (d101, d13, d17);
	nand (d102, d38, d61);
	xnor (d103, d15, d43);
	or (d104, d21, d28);
	and (d105, d34, d66);
	and (d106, d45, d68);
	nand (d107, d19, d63);
	nor (d108, d28, d38);
	and (d109, d14, d23);
	buf (d110, d5);
	not (d111, d21);
	nor (d112, d30, d56);
	xnor (d113, d52, d54);
	buf (d114, d23);
	xnor (d115, d51, d70);
	xor (d116, d36, d67);
	and (d117, d26, d51);
	not (d118, d70);
	nand (d119, d68, d70);
	nand (d120, d18, d65);
	xnor (d121, d62, d69);
	xnor (d122, d27, d33);
	nor (d123, d21, d62);
	xor (d124, d36, d49);
	nor (d125, d26, d53);
	buf (d126, d45);
	and (d127, d17, d36);
	nor (d128, d46, d49);
	buf (d129, d43);
	xnor (d130, d43, d63);
	not (d131, d14);
	nand (d132, d13, d38);
	nand (d133, d12, d60);
	xor (d134, d55, d68);
	buf (d135, d3);
	or (d136, d16, d68);
	nand (d137, d43, d44);
	nor (d138, d55, d64);
	xor (d139, d21, d54);
	and (d140, d36, d57);
	buf (d141, d14);
	xnor (d142, d34, d61);
	nor (d143, d30, d70);
	xor (d144, d56);
	nor (d145, d18, d53);
	xnor (d146, d81, d108);
	xor (d147, d74, d81);
	not (d148, d5);
	xor (d149, d101, d114);
	buf (d150, d112);
	or (d151, d80, d132);
	and (d152, d79, d139);
	or (d153, d82, d142);
	nand (d154, d92, d125);
	nor (d155, d93, d144);
	xor (d156, d90, d132);
	nor (d157, d81, d99);
	not (d158, d138);
	buf (d159, d125);
	or (d160, d97, d115);
	and (d161, d91, d120);
	and (d162, d117, d141);
	and (d163, d102, d106);
	and (d164, d84, d103);
	xnor (d165, d72, d121);
	nor (d166, d106, d129);
	xor (d167, d71, d79);
	and (d168, d126, d144);
	nand (d169, d102, d107);
	nand (d170, d122, d139);
	not (d171, d55);
	and (d172, d115, d127);
	nand (d173, d106, d112);
	or (d174, d90, d126);
	nand (d175, d96, d122);
	xnor (d176, d91, d125);
	nand (d177, d79, d89);
	not (d178, d100);
	or (d179, d76, d115);
	or (d180, d85, d138);
	nand (d181, d91, d111);
	xor (d182, d109, d129);
	buf (d183, d77);
	and (d184, d83, d98);
	nand (d185, d93, d111);
	xor (d186, d109, d145);
	not (d187, d143);
	and (d188, d103, d109);
	nor (d189, d92, d127);
	or (d190, d93, d114);
	not (d191, d26);
	xnor (d192, d74, d141);
	nand (d193, d86, d121);
	buf (d194, d121);
	not (d195, d31);
	buf (d196, d128);
	nand (d197, d75, d96);
	xor (d198, d80, d139);
	xor (d199, d107, d117);
	xor (d200, d129, d133);
	nand (d201, d114, d138);
	xor (d202, d80, d128);
	xor (d203, d89, d143);
	nor (d204, d99, d120);
	nor (d205, d73, d143);
	and (d206, d78, d81);
	buf (d207, d118);
	and (d208, d184, d186);
	not (d209, d107);
	or (d210, d149, d206);
	and (d211, d179, d200);
	or (d212, d163, d207);
	nor (d213, d147, d174);
	buf (d214, d38);
	not (d215, d118);
	xor (d216, d147, d154);
	xor (d217, d163, d206);
	or (d218, d184, d207);
	buf (d219, d18);
	and (d220, d155, d199);
	or (d221, d152, d186);
	xnor (d222, d157, d189);
	not (d223, d65);
	nor (d224, d213, d223);
	and (d225, d214, d221);
	and (d226, d209, d220);
	or (d227, d214, d219);
	nor (d228, d208, d216);
	and (d229, d219, d221);
	buf (d230, d51);
	nor (d231, d215, d220);
	buf (d232, d219);
	buf (d233, d20);
	buf (d234, d110);
	xor (d235, d208, d217);
	buf (d236, d52);
	or (d237, d215, d220);
	xor (d238, d208, d221);
	nor (d239, d212, d222);
	nor (d240, d219, d222);
	xor (d241, d213, d223);
	nor (d242, d208, d223);
	or (d243, d226, d239);
	xnor (d244, d234, d241);
	or (d245, d230, d233);
	nor (d246, d228, d239);
	nand (d247, d231, d236);
	and (d248, d227, d239);
	and (d249, d229, d234);
	xor (d250, d230, d236);
	xnor (d251, d227, d236);
	buf (d252, d28);
	nor (d253, d227, d241);
	nand (d254, d224, d231);
	not (d255, d223);
	not (d256, d212);
	xor (d257, d224, d234);
	buf (d258, d91);
	xnor (d259, d233, d242);
	nor (d260, d227, d229);
	nor (d261, d231, d241);
	or (d262, d226, d234);
	buf (d263, d159);
	buf (d264, d203);
	and (d265, d233, d237);
	nor (d266, d228, d229);
	xor (d267, d233, d236);
	nor (d268, d228, d234);
	and (d269, d230, d236);
	buf (d270, d92);
	xor (d271, d231, d237);
	nor (d272, d226, d227);
	and (d273, d224, d237);
	or (d274, d238, d242);
	and (d275, d228, d237);
	nand (d276, d225, d236);
	nand (d277, d229, d237);
	xor (d278, d224, d241);
	not (d279, d47);
	xnor (d280, d235, d236);
	not (d281, d164);
	xnor (d282, d231, d232);
	xor (d283, d240);
	not (d284, d174);
	not (d285, d120);
	nand (d286, d238, d240);
	nor (d287, d237, d240);
	or (d288, d236, d240);
	nand (d289, d236, d240);
	or (d290, d224, d240);
	buf (d291, d120);
	and (d292, d225, d239);
	xnor (d293, d231);
	xnor (d294, d224, d231);
	nor (d295, d231, d239);
	nand (d296, d232, d236);
	nand (d297, d229, d235);
	not (d298, d114);
	not (d299, d182);
	assign f1 = d297;
	assign f2 = d289;
	assign f3 = d297;
	assign f4 = d299;
	assign f5 = d277;
	assign f6 = d243;
	assign f7 = d286;
	assign f8 = d256;
	assign f9 = d288;
	assign f10 = d283;
endmodule
