module CCGRCG394( x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17, f18, f19, f20, f21, f22, f23, f24, f25, f26 );

	input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17, f18, f19, f20, f21, f22, f23, f24, f25, f26;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314, d315, d316, d317, d318, d319, d320, d321, d322, d323, d324, d325, d326, d327, d328, d329, d330, d331, d332, d333, d334, d335, d336, d337, d338, d339, d340, d341, d342, d343, d344, d345, d346, d347, d348, d349, d350, d351, d352, d353, d354, d355, d356, d357, d358, d359, d360, d361, d362, d363, d364, d365, d366, d367, d368, d369, d370, d371, d372, d373, d374, d375, d376, d377, d378, d379, d380, d381, d382, d383, d384, d385, d386, d387, d388, d389, d390, d391, d392, d393, d394, d395, d396, d397, d398, d399, d400, d401, d402, d403, d404, d405, d406, d407, d408, d409, d410, d411, d412, d413, d414, d415, d416, d417, d418, d419, d420, d421, d422, d423, d424, d425, d426, d427, d428, d429, d430, d431, d432, d433, d434, d435, d436, d437, d438, d439, d440, d441, d442, d443, d444, d445, d446, d447, d448, d449, d450, d451, d452, d453, d454, d455, d456, d457, d458, d459, d460, d461, d462, d463, d464, d465, d466, d467, d468, d469, d470, d471, d472, d473, d474, d475, d476, d477, d478, d479, d480, d481, d482, d483, d484, d485, d486, d487, d488, d489, d490, d491, d492, d493, d494, d495, d496, d497, d498, d499, d500, d501, d502, d503, d504, d505, d506, d507, d508, d509, d510, d511, d512, d513, d514, d515, d516, d517, d518, d519, d520, d521, d522, d523, d524, d525, d526, d527, d528, d529, d530, d531, d532, d533, d534, d535, d536, d537, d538, d539, d540, d541, d542, d543, d544, d545, d546, d547, d548, d549, d550, d551, d552, d553, d554, d555, d556, d557, d558, d559, d560, d561, d562, d563, d564, d565, d566, d567, d568, d569, d570, d571, d572, d573, d574, d575, d576, d577, d578, d579, d580, d581, d582, d583, d584, d585, d586, d587, d588, d589, d590, d591, d592, d593, d594, d595, d596, d597, d598, d599, d600, d601, d602, d603, d604, d605, d606, d607, d608, d609, d610, d611, d612, d613, d614, d615, d616, d617, d618, d619, d620, d621, d622, d623, d624, d625, d626, d627, d628, d629, d630, d631, d632, d633, d634, d635, d636, d637, d638, d639, d640, d641, d642, d643, d644, d645, d646, d647, d648, d649, d650, d651, d652, d653, d654, d655, d656, d657, d658, d659, d660, d661, d662, d663, d664, d665, d666, d667, d668, d669, d670, d671, d672, d673, d674, d675, d676, d677, d678, d679, d680, d681, d682, d683, d684, d685, d686, d687, d688, d689, d690, d691, d692, d693, d694, d695, d696, d697, d698, d699, d700, d701, d702, d703, d704, d705, d706, d707, d708, d709, d710, d711, d712, d713, d714, d715, d716, d717, d718, d719, d720, d721, d722, d723, d724, d725, d726, d727, d728, d729, d730, d731, d732, d733, d734, d735, d736, d737, d738, d739, d740, d741, d742, d743, d744, d745, d746, d747, d748, d749, d750, d751, d752, d753, d754, d755, d756, d757, d758, d759, d760, d761, d762, d763, d764;

	nand ( d1, x1, x13);
	not ( d2, x0);
	and ( d3, x10, x25);
	and ( d4, x1, x16);
	buf ( d5, x4);
	nor ( d6, x16, x26);
	xnor ( d7, x14, x24);
	xor ( d8, x7, x25);
	nor ( d9, x18, x21);
	or ( d10, x14, x27);
	or ( d11, x13, x17);
	and ( d12, x8, x27);
	nor ( d13, x17, x18);
	xnor ( d14, x7, x16);
	nor ( d15, x18, x19);
	not ( d16, x10);
	nand ( d17, x16, x26);
	buf ( d18, x27);
	xnor ( d19, x1, x3);
	not ( d20, x6);
	nand ( d21, x14, x22);
	buf ( d22, x22);
	xnor ( d23, x7, x21);
	xor ( d24, x15, x25);
	or ( d25, x17, x24);
	nor ( d26, x16, x19);
	not ( d27, x26);
	or ( d28, x7, x22);
	xnor ( d29, x3, x13);
	not ( d30, x14);
	or ( d31, x12, x25);
	xor ( d32, x26, x27);
	nor ( d33, x7, x16);
	xor ( d34, x4, x25);
	not ( d35, x18);
	and ( d36, x20, x27);
	buf ( d37, x15);
	nor ( d38, x5, x11);
	not ( d39, x27);
	nor ( d40, x0, x25);
	or ( d41, x6, x22);
	nand ( d42, x17, x23);
	or ( d43, x9, x19);
	nor ( d44, x20, x25);
	or ( d45, x23, x24);
	xor ( d46, x20);
	xnor ( d47, x10, x12);
	nand ( d48, x0, x17);
	or ( d49, x6, x10);
	or ( d50, x0, x10);
	and ( d51, x12, x23);
	and ( d52, x12, x27);
	and ( d53, x18);
	nand ( d54, x10, x26);
	xor ( d55, x0, x4);
	not ( d56, x15);
	or ( d57, x4, x22);
	and ( d58, x1, x11);
	nand ( d59, x9, x27);
	xor ( d60, x11, x14);
	nor ( d61, x1, x3);
	nand ( d62, x17, x27);
	or ( d63, x13, x14);
	buf ( d64, x19);
	buf ( d65, x20);
	and ( d66, x2, x15);
	nor ( d67, x9, x13);
	xor ( d68, d8, d56);
	xor ( d69, d6, d27);
	buf ( d70, x14);
	nand ( d71, d42, d64);
	xor ( d72, d31, d51);
	xor ( d73, d2, d65);
	and ( d74, d11, d31);
	xnor ( d75, d36);
	xor ( d76, d23, d48);
	xor ( d77, d59, d65);
	xnor ( d78, d4, d6);
	buf ( d79, x18);
	nor ( d80, d47, d63);
	xnor ( d81, d3, d24);
	buf ( d82, d42);
	nand ( d83, d28, d36);
	xor ( d84, d4, d20);
	or ( d85, d21, d22);
	xnor ( d86, d53, d59);
	or ( d87, d23, d37);
	xor ( d88, d25, d40);
	xor ( d89, d4, d46);
	xor ( d90, d3, d48);
	nor ( d91, d11, d50);
	not ( d92, d21);
	xor ( d93, d20, d58);
	or ( d94, d16, d47);
	nand ( d95, d15, d43);
	nand ( d96, d24, d64);
	and ( d97, d5, d16);
	and ( d98, d17, d29);
	buf ( d99, d2);
	xnor ( d100, d19, d41);
	not ( d101, x4);
	xnor ( d102, d16, d66);
	nand ( d103, d17, d56);
	and ( d104, d57, d59);
	nand ( d105, d21, d50);
	not ( d106, d7);
	xor ( d107, d4, d10);
	nand ( d108, d55, d60);
	not ( d109, d30);
	and ( d110, d1, d58);
	xor ( d111, d1, d63);
	nand ( d112, d38, d40);
	xor ( d113, d61, d65);
	or ( d114, d23, d25);
	buf ( d115, d13);
	buf ( d116, d9);
	xor ( d117, d52, d63);
	buf ( d118, d51);
	or ( d119, d32, d65);
	or ( d120, d25, d46);
	nand ( d121, d16, d39);
	xor ( d122, d1, d40);
	xnor ( d123, d28, d50);
	nand ( d124, d57, d60);
	nand ( d125, d4, d57);
	and ( d126, d113, d116);
	and ( d127, d72, d103);
	nand ( d128, d80, d98);
	nor ( d129, d92, d102);
	and ( d130, d98, d103);
	or ( d131, d82, d100);
	not ( d132, d25);
	nor ( d133, d83, d120);
	nand ( d134, d105, d112);
	xnor ( d135, d79, d108);
	buf ( d136, d77);
	not ( d137, d37);
	nand ( d138, d98, d115);
	buf ( d139, d3);
	xor ( d140, d73, d108);
	xnor ( d141, d68, d80);
	buf ( d142, d124);
	nor ( d143, d76, d122);
	xor ( d144, d70, d117);
	nand ( d145, d101, d111);
	nor ( d146, d118, d125);
	or ( d147, d97, d103);
	and ( d148, d97, d110);
	nor ( d149, d73, d79);
	xor ( d150, d79, d113);
	buf ( d151, x6);
	nor ( d152, d96, d117);
	and ( d153, d70, d86);
	xor ( d154, d90, d99);
	and ( d155, d85, d90);
	and ( d156, d68, d75);
	or ( d157, d71, d84);
	not ( d158, d79);
	xor ( d159, d69, d83);
	nor ( d160, d78, d80);
	nand ( d161, d68, d74);
	xnor ( d162, d88, d121);
	not ( d163, d110);
	xnor ( d164, d77, d85);
	nand ( d165, d88, d111);
	xor ( d166, d82, d108);
	xor ( d167, d84, d112);
	nor ( d168, d72, d98);
	xnor ( d169, d73, d110);
	or ( d170, d73, d121);
	xor ( d171, d88, d99);
	xor ( d172, d71, d112);
	or ( d173, d115, d122);
	or ( d174, d81, d113);
	nand ( d175, d93, d101);
	xnor ( d176, d80, d82);
	nor ( d177, d73, d107);
	and ( d178, d84, d118);
	xnor ( d179, d111, d115);
	not ( d180, d55);
	xnor ( d181, d75, d119);
	xnor ( d182, d74, d100);
	xnor ( d183, d68, d114);
	nor ( d184, d93, d106);
	nand ( d185, d94, d96);
	or ( d186, d88, d105);
	and ( d187, d72);
	not ( d188, d19);
	and ( d189, d167, d187);
	not ( d190, d177);
	nand ( d191, d142, d173);
	or ( d192, d176, d180);
	xor ( d193, d146, d182);
	not ( d194, d89);
	nor ( d195, d182, d183);
	not ( d196, d156);
	not ( d197, d33);
	or ( d198, d176, d185);
	nand ( d199, d129, d164);
	xnor ( d200, d139, d178);
	xor ( d201, d178, d184);
	xor ( d202, d138, d165);
	and ( d203, d147, d168);
	buf ( d204, d137);
	xnor ( d205, d131, d180);
	not ( d206, x19);
	nand ( d207, d151, d169);
	nor ( d208, d154, d165);
	xnor ( d209, d136, d172);
	nand ( d210, d157, d178);
	xnor ( d211, d172, d177);
	xnor ( d212, d167, d172);
	or ( d213, d163, d169);
	nand ( d214, d144);
	nand ( d215, d166, d176);
	nand ( d216, d190, d204);
	and ( d217, d190, d206);
	xnor ( d218, d199, d209);
	buf ( d219, d17);
	xor ( d220, d189, d212);
	xnor ( d221, d197, d206);
	or ( d222, d193, d197);
	nand ( d223, d189, d197);
	xor ( d224, d198, d207);
	buf ( d225, d86);
	nand ( d226, d199);
	or ( d227, d192, d196);
	or ( d228, d198, d202);
	xor ( d229, d198, d212);
	and ( d230, d197, d205);
	xor ( d231, d189, d202);
	and ( d232, d188, d197);
	not ( d233, x16);
	nand ( d234, d191, d192);
	and ( d235, d189, d209);
	and ( d236, d200, d209);
	not ( d237, x3);
	and ( d238, d188, d206);
	xor ( d239, d194, d212);
	xnor ( d240, d194, d198);
	xor ( d241, d204, d209);
	nand ( d242, d196, d206);
	and ( d243, d189, d208);
	nor ( d244, d202, d210);
	xnor ( d245, d193, d197);
	and ( d246, d192, d206);
	buf ( d247, d5);
	or ( d248, d202, d209);
	nor ( d249, d194, d203);
	and ( d250, d188, d200);
	xnor ( d251, d210, d214);
	or ( d252, d191, d192);
	and ( d253, d202, d203);
	nand ( d254, d199, d203);
	buf ( d255, d186);
	not ( d256, d42);
	xnor ( d257, d197, d201);
	not ( d258, d167);
	buf ( d259, d173);
	or ( d260, d199, d205);
	or ( d261, d197, d215);
	xnor ( d262, d192, d207);
	xnor ( d263, d205, d215);
	buf ( d264, d211);
	and ( d265, d198, d201);
	nor ( d266, d196, d204);
	buf ( d267, d32);
	and ( d268, d189, d200);
	buf ( d269, d177);
	buf ( d270, d190);
	and ( d271, d191, d209);
	or ( d272, d199, d212);
	buf ( d273, d151);
	buf ( d274, d195);
	xor ( d275, d189, d201);
	xnor ( d276, d191, d214);
	nor ( d277, d193, d215);
	nand ( d278, d205, d212);
	nor ( d279, d196, d198);
	xor ( d280, d201, d214);
	not ( d281, d53);
	and ( d282, d201, d202);
	nand ( d283, d232, d265);
	and ( d284, d233, d259);
	nor ( d285, d216, d270);
	buf ( d286, d222);
	or ( d287, d225, d239);
	not ( d288, x9);
	xor ( d289, d262, d268);
	xor ( d290, d254, d268);
	and ( d291, d229, d270);
	xnor ( d292, d233, d236);
	nor ( d293, d228, d265);
	buf ( d294, d215);
	nor ( d295, d219, d231);
	nor ( d296, d225, d271);
	or ( d297, d229, d239);
	nor ( d298, d226, d265);
	or ( d299, d262, d274);
	nand ( d300, d226, d247);
	buf ( d301, d274);
	xor ( d302, d225, d256);
	buf ( d303, d61);
	or ( d304, d245, d263);
	nor ( d305, d220, d244);
	nand ( d306, d249, d258);
	nand ( d307, d217, d277);
	nand ( d308, d240, d244);
	xnor ( d309, d235, d269);
	nor ( d310, d218, d225);
	nand ( d311, d245, d260);
	or ( d312, d237, d275);
	nor ( d313, d266, d280);
	or ( d314, d231, d257);
	nand ( d315, d235, d240);
	nand ( d316, d273, d276);
	nand ( d317, d251, d277);
	xnor ( d318, d242, d281);
	not ( d319, d237);
	nand ( d320, d223, d261);
	not ( d321, d212);
	xor ( d322, d272, d274);
	nand ( d323, d229, d261);
	xor ( d324, d274, d275);
	not ( d325, d265);
	xnor ( d326, d221, d253);
	nand ( d327, d235, d259);
	nand ( d328, d217, d281);
	xor ( d329, d268, d274);
	nor ( d330, d217, d235);
	xor ( d331, d272, d278);
	and ( d332, d238, d248);
	or ( d333, d269, d276);
	nand ( d334, d231, d272);
	xnor ( d335, d271, d276);
	xor ( d336, d243, d267);
	buf ( d337, d119);
	xor ( d338, d262, d281);
	nand ( d339, d240, d241);
	buf ( d340, d280);
	xor ( d341, d267, d277);
	buf ( d342, d72);
	and ( d343, d245, d259);
	nor ( d344, d236, d270);
	buf ( d345, d144);
	or ( d346, d229, d251);
	xnor ( d347, d290, d330);
	xnor ( d348, d297, d303);
	not ( d349, d170);
	not ( d350, d93);
	not ( d351, x7);
	xnor ( d352, d284, d338);
	xor ( d353, d285, d317);
	xor ( d354, d284, d333);
	xor ( d355, d322, d339);
	xor ( d356, d296, d321);
	nor ( d357, d302, d324);
	xor ( d358, d324, d332);
	buf ( d359, d150);
	not ( d360, d16);
	xnor ( d361, d286);
	and ( d362, d339, d346);
	xor ( d363, d302, d340);
	and ( d364, d286, d294);
	buf ( d365, d287);
	nand ( d366, d283, d337);
	nand ( d367, d291, d328);
	and ( d368, d303, d316);
	or ( d369, d300, d322);
	and ( d370, d295, d343);
	xor ( d371, d312, d327);
	xor ( d372, d294, d305);
	xor ( d373, d284, d334);
	buf ( d374, d132);
	xor ( d375, d329, d332);
	and ( d376, d285, d314);
	nor ( d377, d290, d320);
	xnor ( d378, d305, d342);
	xnor ( d379, d325, d328);
	nor ( d380, d301, d319);
	or ( d381, d304, d316);
	xor ( d382, d314, d343);
	and ( d383, d283, d323);
	not ( d384, d297);
	not ( d385, d34);
	not ( d386, d81);
	nand ( d387, d319);
	xnor ( d388, d298);
	xnor ( d389, d317, d328);
	buf ( d390, d175);
	xnor ( d391, d298, d327);
	buf ( d392, d165);
	not ( d393, d77);
	nor ( d394, d305, d323);
	nand ( d395, d291, d301);
	or ( d396, d391);
	nand ( d397, d348, d353);
	nand ( d398, d348, d355);
	or ( d399, d367, d386);
	xor ( d400, d392, d395);
	not ( d401, d54);
	nand ( d402, d362, d369);
	or ( d403, d348, d356);
	xnor ( d404, d371, d392);
	xnor ( d405, d357, d364);
	or ( d406, d348, d389);
	buf ( d407, d241);
	not ( d408, d17);
	xor ( d409, d350, d374);
	xor ( d410, d391);
	and ( d411, d357, d366);
	xnor ( d412, d352, d372);
	nor ( d413, d357, d368);
	nor ( d414, d377, d393);
	xor ( d415, d379, d389);
	xor ( d416, d348, d351);
	xor ( d417, d366, d377);
	and ( d418, d356, d366);
	nor ( d419, d358, d369);
	not ( d420, d301);
	and ( d421, d376, d383);
	buf ( d422, d24);
	xnor ( d423, d367, d379);
	not ( d424, d71);
	not ( d425, d260);
	and ( d426, d357, d385);
	xor ( d427, d349, d385);
	nor ( d428, d347, d376);
	buf ( d429, d356);
	and ( d430, d360, d364);
	or ( d431, d387, d394);
	nor ( d432, d347, d389);
	and ( d433, d354, d357);
	or ( d434, d393, d395);
	xor ( d435, d349, d393);
	or ( d436, d379);
	or ( d437, d375, d383);
	nor ( d438, d362, d366);
	nor ( d439, d380, d387);
	nand ( d440, d365, d379);
	xor ( d441, d372, d386);
	not ( d442, d357);
	nor ( d443, d378, d393);
	or ( d444, d348, d362);
	nor ( d445, d369, d376);
	and ( d446, d364);
	and ( d447, d363, d381);
	or ( d448, d361, d372);
	or ( d449, d371, d392);
	buf ( d450, d96);
	xor ( d451, d397, d442);
	xor ( d452, d412, d427);
	nand ( d453, d416, d443);
	xnor ( d454, d431, d448);
	nand ( d455, d440, d445);
	not ( d456, d330);
	xor ( d457, d399, d404);
	nand ( d458, d407, d444);
	not ( d459, d206);
	buf ( d460, d146);
	buf ( d461, d273);
	and ( d462, d398, d415);
	xor ( d463, d417, d433);
	nor ( d464, d406, d411);
	and ( d465, d418, d425);
	buf ( d466, d52);
	and ( d467, d442);
	xnor ( d468, d413, d421);
	xnor ( d469, d410, d424);
	and ( d470, d407, d419);
	or ( d471, d402, d426);
	xnor ( d472, d406, d427);
	nand ( d473, d437, d447);
	or ( d474, d424, d429);
	or ( d475, d423, d447);
	nor ( d476, d405, d429);
	or ( d477, d396, d403);
	and ( d478, d398, d400);
	nand ( d479, d401, d441);
	not ( d480, d175);
	buf ( d481, d240);
	or ( d482, d402, d443);
	and ( d483, d407, d433);
	or ( d484, d406, d419);
	buf ( d485, d41);
	nand ( d486, d396, d421);
	buf ( d487, d377);
	xor ( d488, d419, d432);
	xnor ( d489, d408, d444);
	and ( d490, d440, d447);
	not ( d491, d2);
	xnor ( d492, d405, d422);
	buf ( d493, d194);
	nand ( d494, d407, d446);
	nor ( d495, d432, d439);
	and ( d496, d398, d410);
	xnor ( d497, d424, d432);
	xnor ( d498, d438, d443);
	nor ( d499, d399, d421);
	nand ( d500, d396, d398);
	and ( d501, d412, d439);
	and ( d502, d406, d416);
	nand ( d503, d409, d448);
	not ( d504, d342);
	not ( d505, d429);
	or ( d506, d400, d412);
	nand ( d507, d398);
	nor ( d508, d420, d442);
	nand ( d509, d421, d431);
	xnor ( d510, d398, d420);
	xnor ( d511, d413, d419);
	xor ( d512, d429, d444);
	xnor ( d513, d404, d408);
	or ( d514, d404, d420);
	or ( d515, d438, d440);
	and ( d516, d422, d449);
	xor ( d517, d401, d435);
	not ( d518, d46);
	xnor ( d519, d455, d495);
	buf ( d520, d11);
	and ( d521, d472, d473);
	buf ( d522, d336);
	or ( d523, d487, d490);
	and ( d524, d451, d452);
	nor ( d525, d502, d517);
	xor ( d526, d501, d502);
	xnor ( d527, d459, d460);
	nand ( d528, d470, d491);
	and ( d529, d460, d483);
	and ( d530, d457, d515);
	xnor ( d531, d465, d480);
	nand ( d532, d459, d462);
	nor ( d533, d473, d510);
	nand ( d534, d452, d498);
	nand ( d535, d464, d514);
	and ( d536, d481, d483);
	nor ( d537, d499, d515);
	not ( d538, d208);
	xnor ( d539, d460, d478);
	buf ( d540, d111);
	nor ( d541, d457, d513);
	or ( d542, d462, d494);
	nand ( d543, d450, d516);
	xnor ( d544, d474, d517);
	nand ( d545, d460, d478);
	xnor ( d546, d492, d497);
	or ( d547, d502, d515);
	buf ( d548, d246);
	not ( d549, d375);
	xnor ( d550, d465, d478);
	nor ( d551, d451, d497);
	nand ( d552, d487, d497);
	xnor ( d553, d467, d508);
	buf ( d554, d324);
	or ( d555, d492, d506);
	or ( d556, d478, d498);
	xnor ( d557, d460, d492);
	xnor ( d558, d472, d509);
	xnor ( d559, d485, d493);
	not ( d560, d88);
	xnor ( d561, d496, d507);
	or ( d562, d466, d509);
	or ( d563, d479, d510);
	nor ( d564, d466, d491);
	and ( d565, d499, d514);
	and ( d566, d456, d506);
	xor ( d567, d522, d550);
	or ( d568, d565, d566);
	or ( d569, d568);
	xnor ( d570, d567);
	not ( d571, d511);
	buf ( d572, d242);
	xnor ( d573, d568);
	nor ( d574, d568);
	nor ( d575, d567);
	xor ( d576, d567);
	buf ( d577, d18);
	nor ( d578, d572, d576);
	or ( d579, d572, d574);
	buf ( d580, d216);
	xor ( d581, d574, d576);
	xnor ( d582, d570, d574);
	xor ( d583, d570, d571);
	xor ( d584, d571, d576);
	xnor ( d585, d569, d576);
	xnor ( d586, d573, d574);
	or ( d587, d570, d572);
	buf ( d588, d344);
	nor ( d589, d570, d573);
	xor ( d590, d571, d574);
	and ( d591, d569, d571);
	not ( d592, d352);
	not ( d593, d137);
	buf ( d594, d125);
	xor ( d595, d571, d575);
	and ( d596, d569, d576);
	buf ( d597, d16);
	or ( d598, d569, d576);
	nand ( d599, d569, d574);
	not ( d600, d219);
	buf ( d601, d576);
	nor ( d602, d569, d576);
	buf ( d603, d239);
	and ( d604, d570, d571);
	buf ( d605, d210);
	and ( d606, d574, d575);
	nor ( d607, d572, d573);
	xor ( d608, d573, d575);
	nand ( d609, d572);
	nor ( d610, d575, d576);
	xnor ( d611, d570, d574);
	nor ( d612, d570, d574);
	nor ( d613, d572, d574);
	nor ( d614, d571, d574);
	nand ( d615, d569, d573);
	xor ( d616, d573, d575);
	or ( d617, d574, d576);
	buf ( d618, d278);
	or ( d619, d571, d572);
	not ( d620, d214);
	xnor ( d621, d573, d575);
	nor ( d622, d571, d576);
	xnor ( d623, d569, d574);
	xnor ( d624, d569, d571);
	xor ( d625, d571, d575);
	not ( d626, d567);
	nand ( d627, d578, d605);
	and ( d628, d577, d613);
	buf ( d629, d319);
	nand ( d630, d596, d623);
	or ( d631, d587);
	buf ( d632, d587);
	nand ( d633, d596, d622);
	and ( d634, d611, d615);
	buf ( d635, d460);
	xor ( d636, d588, d604);
	and ( d637, d598, d610);
	xor ( d638, d604, d624);
	nor ( d639, d595, d618);
	xor ( d640, d587, d610);
	and ( d641, d595, d607);
	nor ( d642, d597, d603);
	and ( d643, d582, d585);
	or ( d644, d584, d591);
	nor ( d645, d595, d613);
	nand ( d646, d603, d611);
	nand ( d647, d578, d580);
	or ( d648, d584, d589);
	not ( d649, d290);
	nor ( d650, d593, d616);
	xor ( d651, d594, d623);
	xnor ( d652, d582, d625);
	buf ( d653, d308);
	not ( d654, d624);
	xor ( d655, d579, d595);
	and ( d656, d602, d623);
	nand ( d657, d578, d600);
	nor ( d658, d583, d613);
	and ( d659, d587, d625);
	nand ( d660, d584, d622);
	or ( d661, d589, d606);
	or ( d662, d583, d589);
	and ( d663, d580, d605);
	nand ( d664, d578, d613);
	xor ( d665, d595, d602);
	not ( d666, d608);
	or ( d667, d579, d620);
	xor ( d668, d587, d603);
	not ( d669, d339);
	nand ( d670, d610, d616);
	buf ( d671, d547);
	or ( d672, d598, d616);
	or ( d673, d589, d622);
	and ( d674, d587, d605);
	buf ( d675, d21);
	not ( d676, d557);
	xnor ( d677, d586, d614);
	and ( d678, d578, d621);
	nor ( d679, d598, d600);
	nor ( d680, d595, d606);
	nor ( d681, d591, d620);
	nand ( d682, d577, d583);
	and ( d683, d597, d604);
	nor ( d684, d582, d612);
	buf ( d685, d340);
	and ( d686, d606, d613);
	buf ( d687, d330);
	and ( d688, d601);
	or ( d689, d593, d618);
	or ( d690, d582, d616);
	and ( d691, d667, d688);
	xnor ( d692, d626, d675);
	or ( d693, d651, d684);
	nand ( d694, d666, d675);
	not ( d695, d305);
	and ( d696, d636, d650);
	nor ( d697, d642, d659);
	nor ( d698, d658);
	nor ( d699, d645, d681);
	nor ( d700, d635, d673);
	and ( d701, d651, d656);
	not ( d702, d672);
	buf ( d703, d297);
	nand ( d704, d664, d665);
	and ( d705, d653, d680);
	or ( d706, d660, d673);
	or ( d707, d650, d654);
	buf ( d708, x10);
	not ( d709, d520);
	and ( d710, d660, d689);
	xnor ( d711, d678, d688);
	or ( d712, d628, d676);
	buf ( d713, d178);
	buf ( d714, d593);
	not ( d715, d252);
	nor ( d716, d627, d641);
	xnor ( d717, d638, d665);
	nor ( d718, d646, d657);
	nor ( d719, d647, d683);
	nor ( d720, d653, d659);
	nor ( d721, d668, d683);
	nand ( d722, d656, d668);
	not ( d723, d504);
	or ( d724, d641, d668);
	nand ( d725, d647, d689);
	buf ( d726, d139);
	or ( d727, d636, d637);
	or ( d728, d663, d674);
	xor ( d729, d657, d674);
	buf ( d730, d372);
	xor ( d731, d650);
	and ( d732, d655, d683);
	or ( d733, d665, d690);
	and ( d734, d650, d676);
	or ( d735, d672, d683);
	xor ( d736, d693, d696);
	xnor ( d737, d701, d717);
	nor ( d738, d721, d734);
	xnor ( d739, d720, d730);
	nor ( d740, d710, d716);
	nand ( d741, d712, d735);
	and ( d742, d705, d721);
	xor ( d743, d710, d734);
	nor ( d744, d691, d720);
	nor ( d745, d691, d718);
	and ( d746, d693, d711);
	not ( d747, d325);
	buf ( d748, x13);
	not ( d749, d727);
	xnor ( d750, d713, d716);
	nand ( d751, d700, d712);
	xnor ( d752, d703, d707);
	nor ( d753, d704, d718);
	nand ( d754, d710, d719);
	xnor ( d755, d721, d724);
	xnor ( d756, d705, d718);
	or ( d757, d695, d729);
	and ( d758, d692, d727);
	nor ( d759, d693, d705);
	xor ( d760, d694, d700);
	xnor ( d761, d715, d727);
	xor ( d762, d695, d718);
	buf ( d763, d747);
	buf ( d764, d78);
	assign f1 = d764;
	assign f2 = d764;
	assign f3 = d764;
	assign f4 = d764;
	assign f5 = d764;
	assign f6 = d764;
	assign f7 = d764;
	assign f8 = d763;
	assign f9 = d763;
	assign f10 = d763;
	assign f11 = d763;
	assign f12 = d764;
	assign f13 = d763;
	assign f14 = d764;
	assign f15 = d764;
	assign f16 = d763;
	assign f17 = d763;
	assign f18 = d763;
	assign f19 = d763;
	assign f20 = d763;
	assign f21 = d764;
	assign f22 = d764;
	assign f23 = d763;
	assign f24 = d764;
	assign f25 = d763;
	assign f26 = d763;
endmodule
