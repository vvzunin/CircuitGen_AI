module CCGRCG36( x0, x1, x2, f1, f2, f3, f4, f5, f6, f7, f8, f9 );

	input x0, x1, x2;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303;

	nand (d1, x1);
	xnor (d2, x0, x2);
	or (d3, x0, x2);
	or (d4, x0, x1);
	and (d5, x1, x2);
	or (d6, x2);
	buf (d7, x1);
	xnor (d8, d6, d7);
	xnor (d9, d1);
	xor (d10, d2, d6);
	or (d11, d7);
	and (d12, d3);
	xor (d13, d2, d4);
	buf (d14, x0);
	xor (d15, d4, d7);
	nand (d16, d5, d6);
	xnor (d17, d3, d6);
	buf (d18, d6);
	or (d19, d2, d5);
	and (d20, d4);
	not (d21, d4);
	xor (d22, d2, d4);
	not (d23, d7);
	nor (d24, d1, d4);
	not (d25, x1);
	and (d26, d1, d7);
	nor (d27, d4, d7);
	nand (d28, d1);
	or (d29, d2, d3);
	and (d30, d4, d6);
	or (d31, d6);
	buf (d32, x2);
	buf (d33, d1);
	buf (d34, d7);
	xnor (d35, d5, d7);
	xnor (d36, d2, d4);
	not (d37, d5);
	xnor (d38, d4);
	nand (d39, d2, d5);
	and (d40, d6);
	nand (d41, d5, d7);
	not (d42, x2);
	and (d43, d2, d4);
	xnor (d44, d1, d2);
	not (d45, d2);
	xnor (d46, d1, d6);
	nor (d47, d2, d7);
	xor (d48, d1, d4);
	nand (d49, d3, d7);
	or (d50, d2);
	and (d51, d1, d2);
	not (d52, d3);
	nand (d53, d3, d5);
	or (d54, d3, d6);
	or (d55, d1, d2);
	or (d56, d25, d46);
	and (d57, d10, d33);
	and (d58, d33, d49);
	or (d59, d31, d48);
	xor (d60, d18, d42);
	xnor (d61, d30, d54);
	nand (d62, d29, d35);
	xnor (d63, d16, d29);
	not (d64, d13);
	or (d65, d11, d33);
	nand (d66, d25, d40);
	buf (d67, d55);
	nor (d68, d26, d28);
	not (d69, d16);
	and (d70, d16, d46);
	not (d71, d25);
	nand (d72, d63, d69);
	xnor (d73, d57, d68);
	nand (d74, d62);
	xor (d75, d59, d67);
	nand (d76, d66, d67);
	or (d77, d69);
	buf (d78, d10);
	not (d79, d35);
	nand (d80, d56, d70);
	not (d81, d57);
	xnor (d82, d56, d70);
	xor (d83, d60, d62);
	or (d84, d68, d69);
	and (d85, d62, d64);
	nand (d86, d59, d63);
	xnor (d87, d64, d70);
	nand (d88, d63, d67);
	nor (d89, d57, d60);
	and (d90, d60, d69);
	xor (d91, d63, d68);
	nand (d92, d57, d58);
	nor (d93, d64, d70);
	xnor (d94, d56, d60);
	nand (d95, d57, d69);
	nand (d96, d67, d70);
	and (d97, d57, d67);
	xnor (d98, d66);
	xnor (d99, d60, d69);
	xnor (d100, d56, d67);
	not (d101, d21);
	nor (d102, d60, d64);
	xnor (d103, d70);
	or (d104, d60, d70);
	or (d105, d67, d70);
	nor (d106, d61, d65);
	nand (d107, d56, d67);
	or (d108, d57, d61);
	and (d109, d58, d60);
	or (d110, d59, d63);
	nand (d111, d60, d68);
	and (d112, d63, d68);
	buf (d113, d33);
	and (d114, d56, d68);
	or (d115, d62, d63);
	buf (d116, d44);
	buf (d117, d48);
	and (d118, d59, d60);
	and (d119, d67, d69);
	nand (d120, d57, d59);
	buf (d121, d19);
	nor (d122, d56, d64);
	and (d123, d101, d103);
	xnor (d124, d104, d112);
	nand (d125, d94, d100);
	nand (d126, d88, d94);
	not (d127, d36);
	nor (d128, d92, d96);
	or (d129, d74, d102);
	buf (d130, d58);
	nor (d131, d71);
	xnor (d132, d84, d88);
	nand (d133, d92, d104);
	xnor (d134, d72, d108);
	xnor (d135, d93, d100);
	xor (d136, d81, d99);
	nand (d137, d91, d122);
	nor (d138, d79, d106);
	xnor (d139, d84, d90);
	nor (d140, d81, d84);
	buf (d141, d115);
	xnor (d142, d97, d113);
	buf (d143, d13);
	and (d144, d77, d98);
	not (d145, d113);
	or (d146, d85, d111);
	nand (d147, d96, d100);
	and (d148, d74, d80);
	xnor (d149, d82, d94);
	buf (d150, d88);
	xor (d151, d93, d104);
	or (d152, d75, d78);
	or (d153, d85, d122);
	buf (d154, d93);
	xor (d155, d91, d96);
	or (d156, d76, d110);
	and (d157, d74, d76);
	xor (d158, d94, d114);
	nand (d159, d98, d100);
	xnor (d160, d102, d115);
	buf (d161, d32);
	nor (d162, d79, d90);
	xnor (d163, d102, d115);
	or (d164, d82, d120);
	xnor (d165, d112, d122);
	or (d166, d102, d115);
	nor (d167, d74, d112);
	nand (d168, d83, d118);
	not (d169, d39);
	nor (d170, d72, d111);
	nand (d171, d78, d108);
	and (d172, d81, d99);
	xor (d173, d79, d92);
	xor (d174, d82, d97);
	buf (d175, d95);
	not (d176, d118);
	and (d177, d80, d111);
	buf (d178, d91);
	and (d179, d101, d117);
	and (d180, d90, d118);
	and (d181, d141, d160);
	xnor (d182, d124, d169);
	buf (d183, d111);
	xnor (d184, d131, d159);
	nor (d185, d127, d155);
	xor (d186, d150, d177);
	nand (d187, d169, d178);
	nand (d188, d136, d179);
	xnor (d189, d128, d164);
	xor (d190, d163, d164);
	not (d191, d163);
	xnor (d192, d133, d146);
	xnor (d193, d160, d171);
	nor (d194, d123, d150);
	buf (d195, d124);
	buf (d196, d12);
	nand (d197, d140, d166);
	xnor (d198, d145, d153);
	nand (d199, d169, d173);
	nand (d200, d158, d172);
	xnor (d201, d162, d175);
	nor (d202, d149, d157);
	nand (d203, d132, d167);
	xor (d204, d127, d171);
	nand (d205, d132, d167);
	xnor (d206, d143, d150);
	nand (d207, d138, d165);
	not (d208, d112);
	xor (d209, d130, d168);
	xor (d210, d140, d165);
	nor (d211, d149, d167);
	xnor (d212, d146, d180);
	xor (d213, d176, d179);
	and (d214, d132, d147);
	xor (d215, d151, d164);
	nor (d216, d140, d166);
	buf (d217, d134);
	buf (d218, d152);
	or (d219, d123, d169);
	xor (d220, d159, d171);
	nor (d221, d129, d145);
	or (d222, d134, d162);
	or (d223, d138, d177);
	xnor (d224, d147, d151);
	xnor (d225, d153, d165);
	xnor (d226, d130, d139);
	nand (d227, d133, d170);
	or (d228, d162, d169);
	not (d229, d139);
	not (d230, d79);
	nor (d231, d133, d152);
	buf (d232, d51);
	xor (d233, d144, d168);
	not (d234, d26);
	and (d235, d153, d165);
	not (d236, d84);
	xor (d237, d137, d152);
	nand (d238, d136, d162);
	buf (d239, d140);
	nor (d240, d149, d174);
	and (d241, d141, d155);
	nor (d242, d125, d136);
	nand (d243, d123, d126);
	nor (d244, d148, d168);
	not (d245, d44);
	xor (d246, d198, d227);
	buf (d247, d132);
	and (d248, d201, d229);
	xnor (d249, d186, d235);
	not (d250, d187);
	xor (d251, d232, d234);
	and (d252, d198, d239);
	and (d253, d219, d243);
	xor (d254, d197, d235);
	nand (d255, d185, d231);
	and (d256, d205, d231);
	xnor (d257, d211, d216);
	not (d258, d30);
	and (d259, d190, d221);
	not (d260, d32);
	not (d261, d95);
	nor (d262, d183, d225);
	buf (d263, d147);
	nand (d264, d185, d231);
	not (d265, d145);
	xor (d266, d184, d192);
	xor (d267, d204, d214);
	or (d268, d181, d189);
	and (d269, d205, d214);
	buf (d270, d209);
	xor (d271, d181, d235);
	buf (d272, d221);
	buf (d273, d64);
	nor (d274, d188, d198);
	not (d275, d182);
	buf (d276, d215);
	not (d277, d117);
	not (d278, d218);
	buf (d279, d40);
	not (d280, d23);
	buf (d281, d63);
	xnor (d282, d181, d198);
	xor (d283, d234, d243);
	nand (d284, d196, d232);
	not (d285, d212);
	nand (d286, d189, d198);
	not (d287, d47);
	not (d288, d105);
	or (d289, d205, d223);
	or (d290, d196, d241);
	or (d291, d231, d240);
	xor (d292, d220, d242);
	or (d293, d231, d243);
	xor (d294, d185, d201);
	buf (d295, d189);
	nor (d296, d195, d225);
	xor (d297, d224, d237);
	and (d298, d224, d231);
	or (d299, d206, d241);
	nor (d300, d219, d230);
	nor (d301, d207, d237);
	or (d302, d192, d215);
	xor (d303, d223, d227);
	assign f1 = d266;
	assign f2 = d248;
	assign f3 = d290;
	assign f4 = d276;
	assign f5 = d299;
	assign f6 = d273;
	assign f7 = d260;
	assign f8 = d290;
	assign f9 = d300;
endmodule
