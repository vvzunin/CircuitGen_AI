module CCGRCG34( x0, x1, x2, f1, f2, f3, f4, f5, f6, f7, f8 );

	input x0, x1, x2;
	output f1, f2, f3, f4, f5, f6, f7, f8;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314, d315, d316, d317, d318, d319, d320, d321, d322, d323, d324, d325, d326, d327, d328, d329, d330, d331, d332, d333, d334, d335, d336, d337, d338, d339, d340, d341, d342, d343, d344, d345, d346, d347, d348, d349, d350, d351, d352, d353, d354, d355, d356, d357, d358, d359, d360, d361, d362, d363, d364, d365, d366, d367, d368, d369, d370, d371, d372, d373, d374, d375, d376, d377, d378, d379, d380, d381, d382, d383, d384, d385;

	buf (d1, x2);
	xnor (d2, x1);
	not (d3, x1);
	buf (d4, x0);
	or (d5, x0, x1);
	nor (d6, x2);
	or (d7, x2);
	nand (d8, x0, x1);
	buf (d9, x1);
	and (d10, x0, x2);
	nand (d11, x2);
	xor (d12, x2);
	xor (d13, x1);
	xor (d14, x0, x2);
	or (d15, x0, x2);
	nor (d16, x1, x2);
	not (d17, x2);
	xor (d18, x0, x1);
	xor (d19, x1, x2);
	and (d20, x1, x2);
	nor (d21, x0, x2);
	or (d22, x1, x2);
	not (d23, d15);
	xor (d24, d15, d21);
	nor (d25, d17, d19);
	and (d26, d7, d10);
	buf (d27, d15);
	or (d28, d8, d14);
	or (d29, d7, d14);
	nor (d30, d13, d22);
	buf (d31, d18);
	xnor (d32, d9, d14);
	xnor (d33, d1, d20);
	nor (d34, d15, d22);
	xnor (d35, d8, d16);
	xnor (d36, d12, d15);
	or (d37, d7, d22);
	nor (d38, d15, d17);
	or (d39, d3, d12);
	xor (d40, d3, d7);
	buf (d41, d14);
	nand (d42, d11, d16);
	not (d43, d19);
	and (d44, d9, d18);
	xor (d45, d7, d19);
	xnor (d46, d5, d10);
	and (d47, d9, d21);
	and (d48, d3, d10);
	and (d49, d11, d21);
	nor (d50, d7, d10);
	nand (d51, d1, d8);
	or (d52, d6, d22);
	not (d53, d2);
	or (d54, d18, d20);
	xor (d55, d10, d18);
	xnor (d56, d4, d10);
	xnor (d57, d15, d16);
	and (d58, d18, d19);
	not (d59, d6);
	and (d60, d8, d15);
	buf (d61, d5);
	nor (d62, d6, d10);
	nand (d63, d2, d18);
	nor (d64, d10, d18);
	or (d65, d12, d15);
	nand (d66, d3, d9);
	xnor (d67, d13, d17);
	not (d68, d1);
	xnor (d69, d1, d19);
	xor (d70, d5, d22);
	xor (d71, d6, d10);
	or (d72, d15, d21);
	nor (d73, d1, d11);
	nand (d74, d13, d20);
	xnor (d75, d15, d19);
	and (d76, d5, d6);
	xnor (d77, d2, d14);
	nand (d78, d17, d22);
	buf (d79, d11);
	nand (d80, d8, d15);
	buf (d81, d16);
	xnor (d82, d2, d17);
	or (d83, d6, d22);
	xnor (d84, d6, d14);
	or (d85, d5, d22);
	xor (d86, d6, d19);
	xor (d87, d9, d20);
	xor (d88, d15, d18);
	nor (d89, d9, d13);
	and (d90, d17, d19);
	xor (d91, d2, d12);
	or (d92, d2, d15);
	xnor (d93, d16, d18);
	xnor (d94, d10, d16);
	xor (d95, d15, d21);
	xnor (d96, d7);
	xnor (d97, d7, d13);
	and (d98, d15, d19);
	nor (d99, d3, d14);
	nor (d100, d7, d19);
	buf (d101, d9);
	nand (d102, d7, d11);
	not (d103, d7);
	nand (d104, d3, d13);
	and (d105, d12, d15);
	xnor (d106, d5, d16);
	not (d107, d91);
	not (d108, d36);
	nand (d109, d57, d66);
	nor (d110, d46, d71);
	or (d111, d29, d54);
	xor (d112, d85, d90);
	xnor (d113, d49, d103);
	nand (d114, d44, d77);
	buf (d115, d87);
	xor (d116, d79, d94);
	nor (d117, d29, d77);
	nand (d118, d28, d90);
	or (d119, d101, d104);
	xor (d120, d27, d85);
	xor (d121, d49, d101);
	not (d122, d75);
	buf (d123, d42);
	and (d124, d111, d113);
	not (d125, d48);
	nor (d126, d107, d115);
	not (d127, d93);
	and (d128, d117, d122);
	and (d129, d110, d116);
	xnor (d130, d113, d115);
	buf (d131, d75);
	or (d132, d115, d122);
	nand (d133, d109, d117);
	not (d134, d106);
	nand (d135, d118, d120);
	or (d136, d111, d115);
	and (d137, d107, d123);
	nand (d138, d112, d115);
	nand (d139, d109, d123);
	or (d140, d117, d120);
	nor (d141, d116, d122);
	xnor (d142, d115, d123);
	xnor (d143, d110, d116);
	or (d144, d110, d119);
	xor (d145, d116);
	nand (d146, d108, d119);
	or (d147, d113, d123);
	not (d148, d64);
	and (d149, d121, d122);
	xnor (d150, d108, d117);
	buf (d151, d69);
	not (d152, d117);
	xnor (d153, d118, d119);
	xnor (d154, d116, d120);
	nor (d155, d107, d114);
	nand (d156, d113, d116);
	buf (d157, d10);
	nor (d158, d115, d123);
	buf (d159, d120);
	xnor (d160, d107, d118);
	and (d161, d117, d123);
	not (d162, d11);
	not (d163, d53);
	xor (d164, d108, d118);
	or (d165, d118, d120);
	xor (d166, d115, d116);
	not (d167, d118);
	nand (d168, d112, d115);
	or (d169, d110, d119);
	or (d170, d108, d117);
	nand (d171, d114, d117);
	xnor (d172, d109, d116);
	buf (d173, d114);
	nand (d174, d108, d112);
	and (d175, d110, d121);
	and (d176, d119, d123);
	or (d177, d110, d111);
	and (d178, d122, d123);
	nor (d179, d111);
	xnor (d180, d109, d112);
	nor (d181, d107, d118);
	not (d182, d62);
	buf (d183, d35);
	nor (d184, d112, d123);
	buf (d185, d103);
	xor (d186, d115, d120);
	xnor (d187, d121, d123);
	xor (d188, d107, d118);
	nand (d189, d107, d120);
	nand (d190, d117, d121);
	xor (d191, d115, d121);
	or (d192, d118, d122);
	buf (d193, d3);
	xnor (d194, d107, d116);
	nor (d195, d117, d121);
	or (d196, d111, d123);
	nor (d197, d109, d110);
	xor (d198, d109, d111);
	not (d199, d25);
	nor (d200, d110, d113);
	nor (d201, d107, d112);
	xnor (d202, d116, d117);
	xnor (d203, d115, d117);
	xor (d204, d116, d119);
	and (d205, d109, d122);
	and (d206, d107, d119);
	xnor (d207, d155, d171);
	buf (d208, d166);
	or (d209, d168, d173);
	xor (d210, d125, d127);
	not (d211, d169);
	not (d212, d28);
	or (d213, d139, d169);
	nor (d214, d156, d177);
	nor (d215, d175, d206);
	nor (d216, d184, d204);
	xor (d217, d186, d189);
	xor (d218, d191, d200);
	nor (d219, d140, d149);
	not (d220, d202);
	buf (d221, d38);
	not (d222, d20);
	nand (d223, d135, d177);
	xor (d224, d170, d194);
	buf (d225, d141);
	nand (d226, d144, d182);
	buf (d227, d107);
	buf (d228, d115);
	nor (d229, d166, d201);
	or (d230, d175, d199);
	or (d231, d164, d205);
	nor (d232, d200, d201);
	nand (d233, d158, d178);
	xnor (d234, d142, d156);
	nand (d235, d136, d150);
	buf (d236, d100);
	nand (d237, d138, d194);
	nor (d238, d136, d161);
	xnor (d239, d210, d222);
	buf (d240, d30);
	nand (d241, d217, d230);
	and (d242, d225, d227);
	nor (d243, d223, d226);
	nand (d244, d221, d230);
	nand (d245, d226, d236);
	buf (d246, d89);
	buf (d247, d90);
	nand (d248, d223, d230);
	xnor (d249, d238);
	nor (d250, d207, d228);
	xor (d251, d231, d236);
	nand (d252, d211, d236);
	xor (d253, d208, d210);
	or (d254, d220, d238);
	nand (d255, d218, d235);
	nand (d256, d221, d231);
	xor (d257, d233, d237);
	nor (d258, d226, d227);
	or (d259, d211, d237);
	buf (d260, d223);
	nor (d261, d211, d236);
	not (d262, d218);
	nand (d263, d209, d230);
	nand (d264, d210, d226);
	nand (d265, d225, d227);
	xor (d266, d208, d225);
	nand (d267, d210, d234);
	nor (d268, d222, d235);
	and (d269, d232, d237);
	buf (d270, d225);
	not (d271, d51);
	nor (d272, d215, d226);
	nand (d273, d217, d222);
	nand (d274, d227, d234);
	xnor (d275, d211, d228);
	nor (d276, d209, d233);
	buf (d277, d179);
	not (d278, d153);
	xor (d279, d223, d234);
	nor (d280, d210, d211);
	nand (d281, d209, d216);
	xor (d282, d211, d232);
	not (d283, d102);
	not (d284, d173);
	or (d285, d218, d227);
	nor (d286, d223, d232);
	buf (d287, d92);
	and (d288, d210, d223);
	xnor (d289, d217, d219);
	xor (d290, d229, d237);
	nor (d291, d208, d225);
	xnor (d292, d223, d227);
	xor (d293, d235, d236);
	nand (d294, d215, d228);
	buf (d295, d113);
	and (d296, d212, d223);
	nand (d297, d223, d236);
	xnor (d298, d226, d236);
	xnor (d299, d217, d226);
	or (d300, d213, d218);
	nor (d301, d221, d226);
	nor (d302, d229, d238);
	xor (d303, d213, d217);
	nand (d304, d208, d231);
	nor (d305, d213, d226);
	xor (d306, d213);
	xnor (d307, d215, d219);
	xnor (d308, d210, d211);
	and (d309, d209, d219);
	and (d310, d209, d215);
	or (d311, d207, d229);
	or (d312, d212, d221);
	or (d313, d220, d238);
	nor (d314, d217, d222);
	xnor (d315, d218, d231);
	or (d316, d207, d216);
	nor (d317, d296, d315);
	xor (d318, d247, d280);
	not (d319, d95);
	buf (d320, d74);
	buf (d321, d227);
	not (d322, d4);
	nand (d323, d259, d291);
	nand (d324, d249, d297);
	not (d325, d297);
	nand (d326, d255, d277);
	nand (d327, d257, d270);
	nand (d328, d277, d305);
	xnor (d329, d279, d313);
	buf (d330, d4);
	or (d331, d273, d314);
	xor (d332, d249, d305);
	xor (d333, d264, d291);
	buf (d334, d158);
	xnor (d335, d255, d299);
	or (d336, d273, d311);
	nand (d337, d290, d303);
	not (d338, d30);
	buf (d339, d66);
	nor (d340, d278, d281);
	xnor (d341, d261, d268);
	not (d342, d292);
	xor (d343, d240, d302);
	not (d344, d32);
	and (d345, d304, d309);
	nor (d346, d246, d288);
	or (d347, d285, d299);
	buf (d348, d277);
	buf (d349, d288);
	nor (d350, d241, d307);
	not (d351, d225);
	or (d352, d251, d310);
	nand (d353, d256, d288);
	buf (d354, d12);
	and (d355, d252, d285);
	nor (d356, d243, d298);
	and (d357, d254, d255);
	buf (d358, d143);
	nor (d359, d272, d275);
	xor (d360, d266, d303);
	buf (d361, d285);
	and (d362, d239, d248);
	xnor (d363, d287, d310);
	not (d364, d165);
	xor (d365, d241, d262);
	buf (d366, d8);
	nor (d367, d291, d311);
	or (d368, d243, d286);
	xnor (d369, d242, d260);
	nand (d370, d267, d299);
	buf (d371, d244);
	nand (d372, d265, d272);
	nor (d373, d252, d295);
	xor (d374, d252, d302);
	xor (d375, d279, d295);
	xnor (d376, d278, d311);
	xor (d377, d296, d308);
	buf (d378, d299);
	xnor (d379, d258, d268);
	nand (d380, d251, d261);
	xnor (d381, d298, d310);
	nor (d382, d289, d296);
	not (d383, d26);
	xnor (d384, d261, d293);
	and (d385, d243, d313);
	assign f1 = d363;
	assign f2 = d325;
	assign f3 = d371;
	assign f4 = d339;
	assign f5 = d379;
	assign f6 = d318;
	assign f7 = d369;
	assign f8 = d328;
endmodule
