module CCGRCG145( x0, x1, x2, x3, x4, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17 );

	input x0, x1, x2, x3, x4;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134;

	buf (d1, x2);
	xor (d2, x3, x4);
	nand (d3, x1, x2);
	xnor (d4, x1, x4);
	not (d5, x2);
	nor (d6, x2);
	nand (d7, x2, x4);
	xnor (d8, x2, x4);
	xor (d9, x2, x3);
	or (d10, x2, x4);
	nand (d11, x0, x3);
	xor (d12, x1, x4);
	and (d13, x1, x3);
	xnor (d14, x0, x1);
	and (d15, x1, x4);
	nand (d16, x0, x1);
	xnor (d17, x0, x3);
	not (d18, x3);
	nand (d19, x0, x2);
	buf (d20, x0);
	xor (d21, x0, x2);
	buf (d22, x3);
	xor (d23, x2, x4);
	nand (d24, x1, x4);
	nand (d25, x0);
	xor (d26, x0, x2);
	or (d27, x3);
	xor (d28, x0, x4);
	or (d29, x0, x1);
	nor (d30, x1);
	not (d31, x4);
	buf (d32, x4);
	and (d33, x0, x1);
	xor (d34, x3, x4);
	nand (d35, x1, x3);
	xor (d36, x1, x3);
	nand (d37, x3);
	xnor (d38, x2, x3);
	xnor (d39, x0, x1);
	or (d40, x1, x2);
	xnor (d41, x3, x4);
	xor (d42, x0, x4);
	nand (d43, x0, x4);
	xnor (d44, x1, x2);
	xor (d45, x0, x3);
	and (d46, x0, x3);
	xnor (d47, x0, x4);
	or (d48, x3, x4);
	or (d49, x0);
	or (d50, x0, x3);
	xnor (d51, d5, d14);
	buf (d52, d25);
	xor (d53, d3, d48);
	buf (d54, d43);
	buf (d55, d34);
	nor (d56, d45, d48);
	nor (d57, d2, d46);
	nand (d58, d3, d13);
	nor (d59, d2, d33);
	or (d60, d15, d22);
	and (d61, d14, d49);
	not (d62, d3);
	nor (d63, d3, d35);
	xnor (d64, d10, d39);
	nor (d65, d1, d10);
	xor (d66, d28, d45);
	nor (d67, d19, d47);
	nor (d68, d22, d30);
	xor (d69, d35, d48);
	not (d70, d21);
	buf (d71, d41);
	xnor (d72, d33, d49);
	nor (d73, d7, d35);
	or (d74, d12, d50);
	nor (d75, d16, d33);
	or (d76, d1, d16);
	nor (d77, d35, d43);
	nand (d78, d11, d42);
	nand (d79, d25, d48);
	xor (d80, d22, d28);
	or (d81, d33, d42);
	nand (d82, d19, d46);
	or (d83, d10, d34);
	or (d84, d35, d36);
	or (d85, d2, d32);
	xnor (d86, d21, d42);
	buf (d87, d74);
	or (d88, d68, d82);
	buf (d89, d49);
	xnor (d90, d64, d75);
	nand (d91, d53, d58);
	buf (d92, d7);
	or (d93, d56, d58);
	nor (d94, d73, d83);
	buf (d95, d16);
	nand (d96, d91, d95);
	nor (d97, d91, d93);
	or (d98, d88, d95);
	not (d99, d23);
	xor (d100, d88, d91);
	nand (d101, d87, d88);
	xnor (d102, d87, d90);
	buf (d103, d14);
	and (d104, d92, d95);
	nor (d105, d91, d92);
	and (d106, d92, d94);
	or (d107, d93);
	not (d108, d62);
	and (d109, d93, d95);
	and (d110, d87, d95);
	nand (d111, d91);
	or (d112, d87, d95);
	or (d113, d94);
	or (d114, d89, d90);
	xnor (d115, d87, d95);
	buf (d116, d20);
	xor (d117, d91, d93);
	not (d118, d15);
	nand (d119, d88, d95);
	nand (d120, d88, d93);
	buf (d121, d19);
	not (d122, d31);
	buf (d123, d13);
	xnor (d124, d89, d95);
	and (d125, d89, d94);
	not (d126, d4);
	buf (d127, d67);
	nor (d128, d92, d95);
	or (d129, d93, d95);
	nand (d130, d91, d95);
	nor (d131, d91, d94);
	or (d132, d89, d92);
	nand (d133, d89, d92);
	not (d134, d12);
	assign f1 = d97;
	assign f2 = d101;
	assign f3 = d97;
	assign f4 = d128;
	assign f5 = d101;
	assign f6 = d113;
	assign f7 = d103;
	assign f8 = d119;
	assign f9 = d116;
	assign f10 = d99;
	assign f11 = d101;
	assign f12 = d122;
	assign f13 = d117;
	assign f14 = d97;
	assign f15 = d128;
	assign f16 = d132;
	assign f17 = d117;
endmodule
