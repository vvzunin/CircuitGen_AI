module CCGRCG153( x0, x1, x2, x3, x4, x5, f1, f2 );

	input x0, x1, x2, x3, x4, x5;
	output f1, f2;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73;

	nor (d1, x0, x4);
	xor (d2, x2, x5);
	and (d3, x0, x3);
	or (d4, x2, x4);
	nor (d5, x5);
	xor (d6, x3);
	buf (d7, x2);
	nor (d8, x3);
	and (d9, x1, x3);
	nand (d10, x0, x2);
	xor (d11, x1, x5);
	not (d12, x2);
	xor (d13, x0, x4);
	xor (d14, x0, x5);
	not (d15, x4);
	or (d16, x2);
	nor (d17, x0, x4);
	nor (d18, x1);
	nor (d19, x1, x5);
	buf (d20, x4);
	xnor (d21, x0, x2);
	and (d22, x1, x2);
	buf (d23, x0);
	nand (d24, x4);
	xor (d25, x0);
	xor (d26, x1, x3);
	or (d27, x0, x4);
	and (d28, x0, x2);
	and (d29, x2, x4);
	buf (d30, x5);
	nand (d31, x1, x2);
	and (d32, x0, x4);
	xor (d33, x1);
	or (d34, x3, x4);
	xor (d35, x0, x3);
	nand (d36, x2, x5);
	xnor (d37, x2, x3);
	xnor (d38, x5);
	buf (d39, x1);
	and (d40, d15, d32);
	not (d41, d21);
	nor (d42, d20, d30);
	buf (d43, d14);
	buf (d44, d3);
	xor (d45, d13, d19);
	nor (d46, d23, d36);
	nor (d47, d4, d14);
	xnor (d48, d34, d35);
	xnor (d49, d32, d36);
	xor (d50, d14, d26);
	buf (d51, d4);
	nor (d52, d31, d36);
	nor (d53, d23, d29);
	or (d54, d21, d30);
	not (d55, d14);
	nand (d56, d6, d24);
	nand (d57, d8, d16);
	nand (d58, d16, d27);
	buf (d59, d17);
	nand (d60, d23, d25);
	and (d61, d27, d34);
	buf (d62, d37);
	nor (d63, d27, d31);
	nand (d64, d8, d39);
	buf (d65, d1);
	or (d66, d18, d23);
	and (d67, d20, d25);
	not (d68, d20);
	or (d69, d28, d34);
	nand (d70, d5, d8);
	nor (d71, d23, d39);
	and (d72, d11, d36);
	and (d73, d3, d24);
	assign f1 = d42;
	assign f2 = d66;
endmodule
