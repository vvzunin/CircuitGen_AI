module CCGRCG21( x0, x1, x2, f1 );

	input x0, x1, x2;
	output f1;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158;

	or (d1, x0);
	xnor (d2, x1);
	and (d3, x1, x2);
	nor (d4, x1);
	nand (d5, x0);
	or (d6, x0, x1);
	nand (d7, x0, x2);
	not (d8, x2);
	and (d9, x1, x2);
	xnor (d10, x0);
	xor (d11, x1, x2);
	nand (d12, x1, x2);
	or (d13, x1, x2);
	xor (d14, x2);
	not (d15, x1);
	nand (d16, x0, x1);
	not (d17, x0);
	xnor (d18, x2);
	nor (d19, x0, x2);
	xnor (d20, x0, x1);
	nand (d21, x1);
	buf (d22, x1);
	buf (d23, x0);
	buf (d24, x2);
	and (d25, x0, x2);
	xor (d26, d2, d18);
	xnor (d27, d1, d18);
	not (d28, d17);
	xor (d29, d2, d6);
	xor (d30, d1, d22);
	nand (d31, d3, d6);
	nand (d32, d4, d15);
	xor (d33, d1, d23);
	nand (d34, d5, d13);
	or (d35, d6, d17);
	xnor (d36, d6);
	nor (d37, d8, d21);
	nand (d38, d3, d24);
	and (d39, d18, d22);
	xor (d40, d2, d24);
	not (d41, d10);
	nand (d42, d13, d19);
	nor (d43, d11, d14);
	buf (d44, d4);
	xor (d45, d14, d24);
	xnor (d46, d4, d22);
	nand (d47, d1, d3);
	and (d48, d10, d13);
	or (d49, d1, d3);
	nor (d50, d7, d25);
	buf (d51, d1);
	nand (d52, d10, d15);
	xnor (d53, d7, d8);
	buf (d54, d18);
	or (d55, d3, d12);
	or (d56, d12, d15);
	nor (d57, d6, d18);
	not (d58, d16);
	xor (d59, d16);
	xor (d60, d9, d20);
	not (d61, d19);
	xnor (d62, d9, d15);
	and (d63, d4, d25);
	xor (d64, d3, d10);
	not (d65, d15);
	not (d66, d2);
	xor (d67, d5, d18);
	and (d68, d15, d20);
	or (d69, d3, d19);
	nor (d70, d7, d8);
	buf (d71, d13);
	nand (d72, d10, d21);
	or (d73, d3, d6);
	nand (d74, d3, d12);
	xor (d75, d11, d19);
	nand (d76, d3, d11);
	nand (d77, d16, d18);
	or (d78, d10, d12);
	not (d79, d20);
	nor (d80, d7, d11);
	not (d81, d22);
	nor (d82, d6, d25);
	nor (d83, d5, d10);
	nor (d84, d2, d4);
	nor (d85, d36, d82);
	xnor (d86, d75, d77);
	xnor (d87, d58, d74);
	xnor (d88, d47, d54);
	nor (d89, d59, d62);
	nor (d90, d82, d83);
	and (d91, d49, d50);
	buf (d92, d44);
	nand (d93, d54, d77);
	xor (d94, d35, d61);
	and (d95, d68, d81);
	buf (d96, d29);
	buf (d97, d75);
	nor (d98, d35, d77);
	nand (d99, d76, d77);
	not (d100, d57);
	nor (d101, d42, d44);
	buf (d102, d27);
	or (d103, d64, d69);
	not (d104, d61);
	nor (d105, d43, d78);
	and (d106, d55, d79);
	or (d107, d46, d63);
	xnor (d108, d41, d59);
	xor (d109, d26, d27);
	xnor (d110, d31, d44);
	buf (d111, d82);
	not (d112, d66);
	not (d113, d25);
	not (d114, d30);
	or (d115, d26, d71);
	not (d116, d39);
	buf (d117, d78);
	buf (d118, d11);
	buf (d119, d66);
	or (d120, d50, d82);
	or (d121, d42, d69);
	nor (d122, d33, d59);
	xnor (d123, d64, d68);
	buf (d124, d37);
	and (d125, d59, d68);
	nor (d126, d79, d84);
	nor (d127, d66, d77);
	xor (d128, d40, d66);
	nand (d129, d49, d55);
	and (d130, d65, d71);
	buf (d131, d80);
	buf (d132, d3);
	and (d133, d41, d64);
	xor (d134, d29, d35);
	not (d135, d55);
	nand (d136, d37, d68);
	xor (d137, d49, d52);
	nand (d138, d26, d54);
	buf (d139, d22);
	buf (d140, d5);
	or (d141, d27, d40);
	xnor (d142, d54, d59);
	nand (d143, d29, d48);
	not (d144, d77);
	xor (d145, d27, d74);
	xor (d146, d63, d74);
	and (d147, d49, d82);
	buf (d148, d40);
	xor (d149, d35, d72);
	buf (d150, d50);
	nand (d151, d39, d83);
	xor (d152, d37, d55);
	xor (d153, d73, d76);
	nand (d154, d45, d68);
	nor (d155, d29, d52);
	and (d156, d49, d78);
	xor (d157, d40, d63);
	xnor (d158, d42, d74);
	assign f1 = d102;
endmodule
