module CCGRCG47( x0, x1, x2, x3, f1, f2, f3, f4 );

	input x0, x1, x2, x3;
	output f1, f2, f3, f4;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240;

	buf (d1, x1);
	xor (d2, x2);
	and (d3, x0, x1);
	nor (d4, x2, x3);
	xnor (d5, x0, x3);
	xnor (d6, x2);
	nor (d7, x3);
	or (d8, x0);
	or (d9, x0, x3);
	xnor (d10, x1, x3);
	nand (d11, x0, x3);
	and (d12, x0, x3);
	xor (d13, x0, x2);
	not (d14, x0);
	nor (d15, x0, x1);
	xor (d16, x0, x1);
	buf (d17, x0);
	nand (d18, x3);
	nand (d19, x0);
	or (d20, x0, x2);
	buf (d21, x2);
	not (d22, x2);
	nand (d23, x2);
	and (d24, x0, x1);
	nand (d25, x1);
	xnor (d26, x0, x2);
	nor (d27, x0, x2);
	nand (d28, x0, x2);
	not (d29, x3);
	or (d30, x1, x2);
	and (d31, x0, x2);
	xor (d32, x3);
	nor (d33, x0, x3);
	xor (d34, x1, x2);
	xnor (d35, x2, x3);
	not (d36, x1);
	or (d37, x1, x2);
	and (d38, x2, x3);
	nand (d39, x0, x1);
	or (d40, x0, x3);
	nor (d41, x1);
	or (d42, x2, x3);
	and (d43, x2, x3);
	and (d44, x1);
	and (d45, d27, d40);
	or (d46, d15, d25);
	xor (d47, d9, d25);
	nor (d48, d13, d38);
	buf (d49, d13);
	nand (d50, d1, d28);
	xor (d51, d2, d30);
	xor (d52, d16, d19);
	or (d53, d14, d18);
	xnor (d54, d31, d37);
	nand (d55, d20, d29);
	xor (d56, d8, d39);
	not (d57, d44);
	xnor (d58, d2, d26);
	nand (d59, d11, d23);
	nor (d60, d11);
	nand (d61, d6, d9);
	nand (d62, d13, d41);
	nor (d63, d9, d19);
	and (d64, d20);
	or (d65, d25, d41);
	and (d66, d5, d28);
	buf (d67, d11);
	xor (d68, d19, d31);
	nor (d69, d17, d43);
	nor (d70, d1, d42);
	nand (d71, d8, d10);
	nand (d72, d11, d36);
	nor (d73, d16, d37);
	buf (d74, d40);
	xor (d75, d10, d27);
	xnor (d76, d6, d8);
	xnor (d77, d38, d42);
	xor (d78, d11, d33);
	xor (d79, d12, d22);
	nand (d80, d13, d44);
	xnor (d81, d39, d40);
	xnor (d82, d11, d31);
	xor (d83, d20, d30);
	xor (d84, d11, d32);
	xnor (d85, d18, d39);
	not (d86, d14);
	nor (d87, d5, d33);
	xor (d88, d2);
	and (d89, d19, d23);
	nand (d90, d27, d28);
	xor (d91, d15, d19);
	or (d92, d23);
	buf (d93, d9);
	xnor (d94, d7, d12);
	or (d95, d17, d36);
	or (d96, d12, d37);
	nor (d97, d39, d41);
	or (d98, d2, d33);
	nand (d99, d17, d19);
	nor (d100, d2, d35);
	xnor (d101, d18, d19);
	not (d102, d99);
	xor (d103, d84, d99);
	nor (d104, d57, d73);
	xor (d105, d51, d55);
	or (d106, d64, d97);
	nor (d107, d70, d99);
	nand (d108, d47, d95);
	not (d109, d71);
	nor (d110, d61, d79);
	nor (d111, d67, d80);
	buf (d112, x3);
	nor (d113, d51, d88);
	or (d114, d70);
	xnor (d115, d63, d89);
	or (d116, d73, d81);
	and (d117, d48, d50);
	or (d118, d55, d64);
	xor (d119, d79, d87);
	xnor (d120, d51, d97);
	xnor (d121, d51, d99);
	or (d122, d65, d82);
	and (d123, d53, d99);
	and (d124, d77, d79);
	buf (d125, d85);
	xor (d126, d90, d99);
	nor (d127, d75, d101);
	or (d128, d75, d87);
	buf (d129, d49);
	xor (d130, d58, d94);
	buf (d131, d39);
	xnor (d132, d65, d70);
	xnor (d133, d50, d100);
	buf (d134, d22);
	nand (d135, d56, d84);
	nand (d136, d59, d81);
	not (d137, d88);
	nand (d138, d46, d82);
	and (d139, d79, d98);
	buf (d140, d70);
	nor (d141, d46, d69);
	and (d142, d62, d64);
	nand (d143, d64, d91);
	xor (d144, d46, d47);
	nor (d145, d46, d74);
	nand (d146, d70, d97);
	nor (d147, d75, d88);
	xor (d148, d73, d81);
	xnor (d149, d84, d99);
	nand (d150, d83, d88);
	buf (d151, d24);
	nor (d152, d72, d93);
	nand (d153, d75, d85);
	or (d154, d59, d63);
	xor (d155, d45, d84);
	or (d156, d88, d99);
	nor (d157, d88, d90);
	not (d158, d75);
	xnor (d159, d49, d93);
	buf (d160, d57);
	nor (d161, d55, d96);
	and (d162, d86, d90);
	xor (d163, d60, d67);
	buf (d164, d45);
	nand (d165, d76, d88);
	nand (d166, d49, d80);
	xnor (d167, d66, d87);
	xor (d168, d84, d101);
	and (d169, d54, d95);
	nand (d170, d73, d82);
	xnor (d171, d123, d145);
	not (d172, d146);
	or (d173, d143, d168);
	nand (d174, d103, d133);
	nor (d175, d116, d168);
	xor (d176, d143, d158);
	buf (d177, d136);
	or (d178, d111, d161);
	or (d179, d115, d158);
	nand (d180, d119, d137);
	and (d181, d116, d154);
	xnor (d182, d114, d120);
	nor (d183, d117, d140);
	nor (d184, d123, d131);
	nor (d185, d119, d142);
	xnor (d186, d166, d169);
	or (d187, d130, d144);
	buf (d188, d83);
	nor (d189, d122, d140);
	xnor (d190, d148, d154);
	not (d191, d86);
	or (d192, d130, d135);
	or (d193, d152, d164);
	xor (d194, d140, d154);
	buf (d195, d30);
	not (d196, d36);
	xnor (d197, d106, d137);
	xor (d198, d102, d161);
	and (d199, d111, d128);
	xnor (d200, d114, d120);
	not (d201, d43);
	buf (d202, d34);
	or (d203, d106, d136);
	xor (d204, d109, d138);
	and (d205, d139, d144);
	and (d206, d116, d136);
	nor (d207, d110, d170);
	buf (d208, d129);
	or (d209, d102, d125);
	or (d210, d102, d116);
	nand (d211, d129, d145);
	xor (d212, d120, d158);
	xnor (d213, d109, d130);
	nor (d214, d122, d136);
	or (d215, d134, d135);
	nor (d216, d118, d163);
	not (d217, d108);
	xnor (d218, d136, d163);
	nor (d219, d126, d146);
	buf (d220, d134);
	nor (d221, d127, d154);
	xor (d222, d112, d150);
	xor (d223, d158, d170);
	nor (d224, d138, d144);
	nor (d225, d131, d167);
	and (d226, d137, d144);
	xor (d227, d140, d144);
	buf (d228, d73);
	or (d229, d137, d149);
	xor (d230, d146, d165);
	nand (d231, d113, d154);
	and (d232, d131, d154);
	or (d233, d104, d137);
	not (d234, d20);
	or (d235, d131, d161);
	not (d236, d151);
	xnor (d237, d157, d164);
	and (d238, d128, d132);
	and (d239, d142, d165);
	not (d240, d119);
	assign f1 = d206;
	assign f2 = d193;
	assign f3 = d232;
	assign f4 = d187;
endmodule
