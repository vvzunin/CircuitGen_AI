module CCGRCG176( x0, x1, x2, x3, x4, x5, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14 );

	input x0, x1, x2, x3, x4, x5;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314, d315, d316, d317, d318, d319, d320, d321, d322, d323, d324, d325, d326, d327, d328, d329, d330, d331, d332, d333, d334, d335, d336, d337, d338, d339, d340, d341, d342, d343, d344, d345, d346, d347, d348, d349, d350, d351, d352, d353, d354, d355, d356, d357, d358, d359, d360, d361, d362, d363, d364, d365, d366, d367, d368, d369, d370, d371, d372, d373, d374, d375, d376, d377, d378, d379, d380, d381;

	nand (d1, x1, x2);
	nor (d2, x2, x3);
	not (d3, x1);
	buf (d4, x3);
	buf (d5, x2);
	nor (d6, x1, x2);
	xor (d7, x0);
	buf (d8, x0);
	and (d9, x0, x1);
	nand (d10, x3, x5);
	and (d11, x0, x2);
	xor (d12, x1, x5);
	nand (d13, x3);
	nor (d14, x2, x4);
	xor (d15, x4, x5);
	nor (d16, x2, x4);
	xor (d17, x1, x2);
	nand (d18, x2, x3);
	buf (d19, x1);
	xnor (d20, x1, x5);
	not (d21, x2);
	xor (d22, x0, x2);
	not (d23, x4);
	xor (d24, x0, x5);
	and (d25, x4, x5);
	xnor (d26, x4, x5);
	nand (d27, x0, x1);
	xnor (d28, x0, x4);
	and (d29, x2, x4);
	nor (d30, x1, x4);
	xnor (d31, x1, x4);
	nor (d32, x2);
	and (d33, x0, x5);
	nor (d34, x1, x5);
	or (d35, x0, x1);
	xnor (d36, x2, x5);
	nor (d37, x1, x3);
	or (d38, x0);
	and (d39, x3);
	xnor (d40, x1, x2);
	or (d41, x2, x4);
	xor (d42, x2);
	xnor (d43, x4, x5);
	not (d44, x3);
	xnor (d45, x2, x4);
	and (d46, x0, x5);
	or (d47, x2, x3);
	or (d48, x1, x2);
	and (d49, x4, x5);
	nand (d50, x0, x5);
	and (d51, x2, x3);
	nand (d52, x1, x4);
	nand (d53, x1, x3);
	and (d54, x3, x4);
	nand (d55, x3, x4);
	not (d56, x5);
	xor (d57, x3, x5);
	nor (d58, x3, x5);
	nand (d59, x0, x5);
	xnor (d60, x3, x5);
	xor (d61, x3);
	nand (d62, x0);
	or (d63, x3, x5);
	nand (d64, x4);
	and (d65, x2, x4);
	xnor (d66, x5);
	not (d67, x0);
	xor (d68, d1, d23);
	buf (d69, d32);
	buf (d70, d17);
	and (d71, d36, d58);
	and (d72, d25, d29);
	not (d73, d29);
	and (d74, d43, d54);
	not (d75, d37);
	not (d76, d28);
	nor (d77, d7, d53);
	or (d78, d17, d54);
	buf (d79, d57);
	xnor (d80, d22, d28);
	nand (d81, d17, d56);
	not (d82, d52);
	not (d83, d2);
	xor (d84, d19, d62);
	not (d85, d44);
	xnor (d86, d42, d58);
	and (d87, d27, d43);
	nand (d88, d16, d63);
	not (d89, d35);
	nor (d90, d35, d40);
	xor (d91, d19, d43);
	and (d92, d6, d10);
	and (d93, d23, d46);
	not (d94, d15);
	nand (d95, d55, d66);
	buf (d96, d23);
	buf (d97, d62);
	not (d98, d60);
	and (d99, d12, d36);
	buf (d100, d15);
	nor (d101, d29, d60);
	and (d102, d4, d30);
	nor (d103, d53, d59);
	nand (d104, d14, d50);
	buf (d105, x4);
	or (d106, d38, d62);
	buf (d107, d58);
	buf (d108, x5);
	nor (d109, d42, d65);
	xor (d110, d8, d29);
	nand (d111, d58, d63);
	xnor (d112, d7, d65);
	xor (d113, d36, d43);
	nor (d114, d13, d28);
	not (d115, d8);
	and (d116, d2, d42);
	nand (d117, d10, d47);
	xnor (d118, d42, d63);
	buf (d119, d55);
	not (d120, d25);
	and (d121, d34, d55);
	or (d122, d10, d51);
	xor (d123, d7, d19);
	and (d124, d18, d40);
	or (d125, d25, d46);
	buf (d126, d35);
	or (d127, d47, d65);
	xnor (d128, d54, d62);
	buf (d129, d24);
	xor (d130, d36, d63);
	xnor (d131, d4, d33);
	xnor (d132, d22, d48);
	xor (d133, d1, d55);
	not (d134, d5);
	nand (d135, d43, d64);
	and (d136, d39, d61);
	xor (d137, d36, d54);
	not (d138, d55);
	or (d139, d30, d57);
	and (d140, d48, d55);
	not (d141, d12);
	nand (d142, d19, d49);
	xor (d143, d22, d52);
	and (d144, d20, d39);
	nand (d145, d17, d47);
	xnor (d146, d8, d36);
	buf (d147, d2);
	buf (d148, d29);
	nor (d149, d36, d52);
	nor (d150, d6, d34);
	nand (d151, d11, d32);
	xor (d152, d31, d45);
	xor (d153, d1, d19);
	buf (d154, d53);
	and (d155, d4, d48);
	and (d156, d5, d17);
	and (d157, d10, d62);
	or (d158, d29, d56);
	or (d159, d23, d65);
	and (d160, d106, d112);
	buf (d161, d127);
	xor (d162, d90, d121);
	nand (d163, d132, d134);
	or (d164, d102, d119);
	and (d165, d79, d91);
	or (d166, d90);
	xnor (d167, d83, d105);
	nor (d168, d96, d99);
	not (d169, d86);
	nand (d170, d69, d76);
	xor (d171, d132, d152);
	buf (d172, d113);
	nor (d173, d83, d88);
	or (d174, d86, d127);
	nor (d175, d106, d137);
	xor (d176, d119, d152);
	nand (d177, d82, d109);
	xor (d178, d68, d69);
	xnor (d179, d72, d101);
	xnor (d180, d147, d158);
	and (d181, d122, d138);
	xnor (d182, d80, d106);
	xor (d183, d92, d134);
	buf (d184, d61);
	nand (d185, d102, d108);
	buf (d186, d14);
	nand (d187, d146, d157);
	not (d188, d89);
	buf (d189, d132);
	xor (d190, d77, d95);
	xnor (d191, d80, d100);
	and (d192, d68, d98);
	or (d193, d134, d155);
	xnor (d194, d92, d100);
	or (d195, d86, d133);
	xor (d196, d73, d79);
	nor (d197, d68, d120);
	nand (d198, d126, d157);
	or (d199, d106, d110);
	nor (d200, d116, d151);
	or (d201, d99, d107);
	not (d202, d103);
	nor (d203, d141, d149);
	buf (d204, d41);
	xnor (d205, d70, d152);
	nand (d206, d70, d133);
	not (d207, d147);
	nand (d208, d70, d112);
	not (d209, d142);
	not (d210, d143);
	and (d211, d107, d147);
	xnor (d212, d90, d134);
	xnor (d213, d134, d158);
	nand (d214, d71, d93);
	nand (d215, d91, d128);
	or (d216, d113, d117);
	xnor (d217, d72, d84);
	xnor (d218, d121, d133);
	not (d219, d106);
	xor (d220, d81, d101);
	xor (d221, d98, d113);
	or (d222, d151, d154);
	buf (d223, d165);
	xnor (d224, d165, d185);
	xor (d225, d163, d174);
	xnor (d226, d163, d186);
	xnor (d227, d185, d217);
	nand (d228, d175, d203);
	nand (d229, d178, d197);
	or (d230, d169, d191);
	xor (d231, d194, d215);
	xnor (d232, d211, d213);
	and (d233, d173, d222);
	or (d234, d204, d205);
	not (d235, d189);
	buf (d236, d56);
	not (d237, d197);
	and (d238, d177, d218);
	and (d239, d161, d174);
	xnor (d240, d200, d215);
	or (d241, d207, d215);
	xor (d242, d165, d205);
	not (d243, d70);
	buf (d244, d39);
	xnor (d245, d203, d213);
	not (d246, d171);
	or (d247, d173, d221);
	xor (d248, d180, d195);
	nor (d249, d211, d219);
	nor (d250, d213, d214);
	nor (d251, d185, d191);
	buf (d252, d52);
	and (d253, d161, d191);
	xor (d254, d168, d177);
	or (d255, d211, d218);
	nor (d256, d204, d213);
	nand (d257, d193, d198);
	nor (d258, d182, d187);
	nand (d259, d181, d192);
	not (d260, d207);
	buf (d261, d44);
	xor (d262, d163, d219);
	nand (d263, d195, d215);
	nand (d264, d160, d184);
	and (d265, d161, d165);
	xnor (d266, d179, d216);
	or (d267, d198, d212);
	nor (d268, d219, d222);
	and (d269, d209, d220);
	and (d270, d188, d189);
	nor (d271, d161, d213);
	xnor (d272, d197, d199);
	xor (d273, d170, d220);
	nor (d274, d161, d199);
	nand (d275, d188, d219);
	or (d276, d169, d194);
	and (d277, d187, d197);
	nor (d278, d167, d202);
	xor (d279, d175, d186);
	nand (d280, d179, d207);
	not (d281, d56);
	not (d282, d135);
	not (d283, d61);
	buf (d284, d8);
	nor (d285, d276, d279);
	xor (d286, d247, d260);
	and (d287, d253, d280);
	buf (d288, d245);
	nor (d289, d246, d272);
	nor (d290, d231, d265);
	xnor (d291, d238, d239);
	or (d292, d246, d249);
	not (d293, d211);
	xor (d294, d239, d241);
	and (d295, d273, d281);
	nand (d296, d232, d271);
	xnor (d297, d245, d253);
	xnor (d298, d266, d277);
	buf (d299, d153);
	xnor (d300, d226, d240);
	nand (d301, d242, d262);
	nor (d302, d266, d267);
	nand (d303, d241, d265);
	xnor (d304, d224, d241);
	or (d305, d230, d244);
	nand (d306, d260, d282);
	buf (d307, d261);
	buf (d308, d94);
	nand (d309, d256, d259);
	and (d310, d262, d276);
	or (d311, d247, d249);
	buf (d312, d240);
	not (d313, d280);
	buf (d314, d75);
	buf (d315, d96);
	and (d316, d243, d262);
	xnor (d317, d225, d255);
	buf (d318, d137);
	nand (d319, d259, d269);
	buf (d320, d233);
	and (d321, d224, d281);
	and (d322, d235, d261);
	not (d323, d205);
	and (d324, d256, d269);
	buf (d325, d10);
	nor (d326, d239, d248);
	not (d327, d203);
	or (d328, d255, d281);
	or (d329, d230, d278);
	nand (d330, d253, d262);
	nor (d331, d274, d278);
	xnor (d332, d229, d252);
	nor (d333, d253, d281);
	nand (d334, d235, d260);
	xnor (d335, d230, d236);
	xnor (d336, d224, d275);
	buf (d337, d241);
	nand (d338, d225, d233);
	xnor (d339, d226, d281);
	not (d340, d228);
	or (d341, d272, d283);
	and (d342, d244, d255);
	and (d343, d245, d255);
	xnor (d344, d237, d240);
	xor (d345, d224, d247);
	xnor (d346, d262, d277);
	nand (d347, d246, d247);
	buf (d348, d59);
	buf (d349, d131);
	xor (d350, d241, d273);
	not (d351, d151);
	not (d352, d100);
	nor (d353, d240, d257);
	nand (d354, d242, d248);
	not (d355, d98);
	xnor (d356, d242, d266);
	buf (d357, d251);
	nor (d358, d224, d282);
	not (d359, d241);
	nand (d360, d248, d277);
	xor (d361, d249, d280);
	xnor (d362, d232, d284);
	and (d363, d227, d270);
	buf (d364, d142);
	or (d365, d245, d255);
	buf (d366, d169);
	nand (d367, d240, d241);
	nor (d368, d239, d249);
	or (d369, d253, d269);
	xnor (d370, d234, d260);
	xor (d371, d246, d270);
	or (d372, d226, d265);
	not (d373, d104);
	xor (d374, d242, d269);
	nand (d375, d233, d278);
	buf (d376, d246);
	nand (d377, d241, d262);
	buf (d378, d97);
	or (d379, d236, d247);
	nand (d380, d242, d272);
	buf (d381, d101);
	assign f1 = d308;
	assign f2 = d366;
	assign f3 = d292;
	assign f4 = d352;
	assign f5 = d354;
	assign f6 = d291;
	assign f7 = d332;
	assign f8 = d362;
	assign f9 = d358;
	assign f10 = d350;
	assign f11 = d365;
	assign f12 = d300;
	assign f13 = d293;
	assign f14 = d299;
endmodule
