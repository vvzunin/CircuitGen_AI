module CCGRCG93( x0, x1, x2, x3, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10 );

	input x0, x1, x2, x3;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314, d315, d316, d317, d318, d319, d320, d321, d322, d323, d324, d325, d326, d327, d328, d329, d330, d331, d332, d333, d334, d335, d336, d337, d338, d339, d340, d341, d342, d343, d344, d345, d346, d347, d348, d349, d350, d351, d352, d353, d354, d355, d356, d357, d358, d359, d360, d361, d362, d363, d364, d365, d366, d367, d368, d369, d370, d371, d372, d373, d374, d375, d376, d377, d378, d379, d380, d381, d382, d383, d384, d385, d386, d387, d388, d389, d390, d391, d392, d393, d394, d395, d396, d397, d398, d399, d400, d401, d402, d403, d404, d405, d406, d407, d408, d409, d410, d411, d412, d413, d414, d415, d416, d417, d418, d419, d420, d421, d422, d423, d424, d425, d426, d427, d428, d429, d430, d431, d432, d433, d434, d435, d436, d437, d438, d439, d440, d441, d442, d443, d444, d445, d446, d447, d448, d449, d450, d451, d452, d453, d454, d455, d456, d457, d458, d459, d460, d461, d462, d463, d464, d465, d466, d467, d468, d469, d470, d471, d472, d473, d474, d475, d476, d477, d478, d479, d480, d481, d482, d483, d484, d485, d486, d487, d488, d489, d490, d491, d492, d493, d494, d495, d496, d497, d498, d499, d500, d501, d502, d503, d504, d505, d506, d507, d508, d509, d510, d511, d512, d513, d514, d515, d516, d517, d518, d519, d520, d521, d522, d523, d524, d525, d526, d527, d528, d529, d530, d531, d532, d533, d534, d535, d536, d537, d538, d539, d540, d541, d542, d543, d544, d545, d546, d547, d548, d549, d550, d551, d552, d553, d554, d555, d556, d557, d558, d559, d560, d561, d562, d563, d564, d565, d566, d567, d568, d569, d570;

	or (d1, x0, x2);
	nor (d2, x0, x3);
	and (d3, x1, x3);
	xnor (d4, x2, x3);
	nand (d5, x0);
	or (d6, x2, x3);
	xnor (d7, x1, x2);
	xor (d8, x0, x2);
	and (d9, x1, x2);
	or (d10, x0, x3);
	xor (d11, x0);
	and (d12, x0, x2);
	nand (d13, x2, x3);
	buf (d14, x0);
	xor (d15, x0, x2);
	nor (d16, x0, x3);
	not (d17, x3);
	and (d18, x3);
	nor (d19, x1, x3);
	and (d20, x0, x3);
	nor (d21, x3);
	or (d22, x1, x3);
	nand (d23, x2);
	not (d24, x2);
	and (d25, x2, x3);
	xor (d26, x0, x3);
	nor (d27, x1);
	or (d28, x2);
	xnor (d29, x0, x3);
	nor (d30, x1, x2);
	xnor (d31, x3);
	buf (d32, x2);
	buf (d33, x3);
	nand (d34, x2, x3);
	nand (d35, x1, x2);
	xnor (d36, x1);
	not (d37, x0);
	nor (d38, x0, x2);
	or (d39, x0);
	nor (d40, x2, x3);
	xor (d41, x1, x3);
	nor (d42, x0, x1);
	xnor (d43, x0, x3);
	nand (d44, x0, x3);
	not (d45, x1);
	nor (d46, x2, x3);
	nand (d47, x0, x2);
	nor (d48, x0);
	xnor (d49, x0, x2);
	or (d50, x1, x3);
	xor (d51, x0, x3);
	nand (d52, x1);
	and (d53, x0, x1);
	xor (d54, x1, x3);
	or (d55, x1, x2);
	nand (d56, x0, x1);
	buf (d57, x1);
	xor (d58, x3);
	or (d59, x2, x3);
	xnor (d60, x1, x3);
	or (d61, x1);
	xnor (d62, x0, x1);
	or (d63, x1, x2);
	and (d64, x1, x3);
	and (d65, x1);
	or (d66, x0, x2);
	buf (d67, d56);
	buf (d68, d61);
	or (d69, d39, d52);
	xor (d70, d7, d10);
	nand (d71, d35, d48);
	nand (d72, d26, d60);
	buf (d73, d11);
	xor (d74, d39, d64);
	buf (d75, d50);
	and (d76, d4, d49);
	and (d77, d18, d52);
	and (d78, d41, d49);
	xor (d79, d8, d30);
	nor (d80, d46, d64);
	or (d81, d28, d49);
	and (d82, d55, d63);
	xnor (d83, d47, d52);
	nand (d84, d17, d54);
	not (d85, d18);
	xor (d86, d21, d31);
	nor (d87, d8, d43);
	or (d88, d24, d39);
	nor (d89, d21, d61);
	xor (d90, d33, d36);
	xor (d91, d3, d41);
	and (d92, d16, d51);
	and (d93, d10, d49);
	and (d94, d9, d43);
	xor (d95, d10, d36);
	and (d96, d17, d28);
	xor (d97, d6, d12);
	nor (d98, d22, d36);
	and (d99, d1, d39);
	buf (d100, d65);
	and (d101, d26, d47);
	xor (d102, d46, d53);
	xor (d103, d6, d34);
	not (d104, d19);
	buf (d105, d5);
	and (d106, d3, d5);
	buf (d107, d45);
	and (d108, d11, d51);
	buf (d109, d18);
	nor (d110, d16, d49);
	and (d111, d41, d42);
	nor (d112, d3, d29);
	nand (d113, d12, d47);
	buf (d114, d49);
	not (d115, d7);
	not (d116, d17);
	not (d117, d3);
	nand (d118, d1, d28);
	and (d119, d36, d63);
	nor (d120, d42, d53);
	xor (d121, d37, d48);
	or (d122, d25, d58);
	xor (d123, d37, d66);
	not (d124, d63);
	buf (d125, d53);
	not (d126, d25);
	or (d127, d9, d39);
	nor (d128, d26, d52);
	or (d129, d37, d41);
	nand (d130, d9, d27);
	nor (d131, d10, d47);
	nand (d132, d86, d110);
	or (d133, d72, d75);
	or (d134, d108, d112);
	not (d135, d62);
	buf (d136, d38);
	nand (d137, d82, d113);
	xnor (d138, d92, d95);
	and (d139, d80, d109);
	nand (d140, d95, d108);
	and (d141, d112, d127);
	and (d142, d119, d124);
	nor (d143, d81, d100);
	xnor (d144, d74, d113);
	buf (d145, d19);
	not (d146, d125);
	or (d147, d104, d120);
	or (d148, d123, d125);
	buf (d149, d101);
	and (d150, d72, d106);
	nand (d151, d67, d115);
	or (d152, d96, d107);
	nor (d153, d100, d112);
	and (d154, d87, d128);
	not (d155, d39);
	nor (d156, d96, d110);
	and (d157, d105, d125);
	buf (d158, d28);
	nand (d159, d126, d129);
	xor (d160, d79, d115);
	nor (d161, d70, d115);
	xor (d162, d107, d119);
	xnor (d163, d78, d112);
	nor (d164, d75, d128);
	and (d165, d102, d112);
	xor (d166, d85, d115);
	nand (d167, d75, d80);
	or (d168, d87, d103);
	xor (d169, d88, d109);
	nor (d170, d116, d125);
	not (d171, d33);
	nor (d172, d75, d79);
	and (d173, d87, d125);
	and (d174, d73, d98);
	nand (d175, d84, d93);
	and (d176, d97, d114);
	not (d177, d4);
	nor (d178, d68);
	and (d179, d95);
	and (d180, d114, d128);
	xnor (d181, d92, d93);
	or (d182, d97, d108);
	not (d183, d73);
	buf (d184, d114);
	not (d185, d2);
	buf (d186, d27);
	buf (d187, d123);
	nor (d188, d114, d119);
	xnor (d189, d75, d121);
	nand (d190, d124, d131);
	or (d191, d83, d116);
	and (d192, d89, d129);
	not (d193, d29);
	and (d194, d99, d122);
	and (d195, d110, d125);
	nor (d196, d86, d91);
	or (d197, d71);
	or (d198, d111, d130);
	xnor (d199, d70, d125);
	and (d200, d85, d95);
	and (d201, d96, d113);
	nand (d202, d87, d88);
	buf (d203, d44);
	nor (d204, d91, d109);
	xor (d205, d71, d113);
	nand (d206, d105, d113);
	nor (d207, d96, d106);
	and (d208, d79, d125);
	nand (d209, d156, d168);
	not (d210, d202);
	xnor (d211, d142, d164);
	xnor (d212, d180, d189);
	nor (d213, d136, d165);
	xor (d214, d188, d199);
	xnor (d215, d181, d184);
	not (d216, d138);
	nand (d217, d166, d204);
	xor (d218, d157, d162);
	not (d219, d98);
	not (d220, d21);
	xor (d221, d161, d191);
	xor (d222, d141, d142);
	and (d223, d185, d204);
	nor (d224, d155, d203);
	nor (d225, d184, d203);
	xnor (d226, d144, d199);
	xnor (d227, d136, d149);
	xnor (d228, d189, d196);
	xnor (d229, d139, d187);
	xor (d230, d153, d180);
	nand (d231, d193, d197);
	nor (d232, d198, d205);
	buf (d233, d122);
	not (d234, d59);
	nand (d235, d171, d199);
	xnor (d236, d135, d136);
	xnor (d237, d167, d197);
	xor (d238, d175, d176);
	xnor (d239, d195, d196);
	not (d240, d44);
	or (d241, d146, d190);
	not (d242, d191);
	and (d243, d179, d187);
	and (d244, d135, d147);
	nor (d245, d194, d199);
	or (d246, d158, d187);
	or (d247, d169, d186);
	nor (d248, d148, d180);
	not (d249, d161);
	buf (d250, d78);
	buf (d251, d115);
	nand (d252, d145);
	not (d253, d61);
	and (d254, d150, d192);
	xnor (d255, d156, d205);
	not (d256, d76);
	xnor (d257, d217, d254);
	xnor (d258, d214, d253);
	or (d259, d214, d244);
	xor (d260, d243, d253);
	nand (d261, d226, d254);
	and (d262, d222, d229);
	or (d263, d220, d247);
	and (d264, d242, d247);
	or (d265, d229, d242);
	nand (d266, d232, d241);
	nor (d267, d215, d225);
	xnor (d268, d250, d253);
	nand (d269, d221, d225);
	buf (d270, d29);
	xnor (d271, d240, d245);
	or (d272, d218, d235);
	buf (d273, d68);
	not (d274, d47);
	xnor (d275, d225, d249);
	or (d276, d232, d246);
	nand (d277, d221, d226);
	xnor (d278, d228, d250);
	and (d279, d233, d234);
	xnor (d280, d214, d232);
	and (d281, d226, d236);
	and (d282, d224, d228);
	nor (d283, d226, d247);
	and (d284, d224, d241);
	nor (d285, d217, d232);
	xnor (d286, d209, d212);
	nor (d287, d228, d248);
	buf (d288, d238);
	buf (d289, d193);
	nand (d290, d210, d228);
	nand (d291, d220, d253);
	xnor (d292, d242, d250);
	nor (d293, d222, d247);
	xor (d294, d238, d249);
	xor (d295, d228, d250);
	not (d296, d181);
	nor (d297, d228, d252);
	nor (d298, d213, d222);
	or (d299, d222, d241);
	and (d300, d219, d244);
	buf (d301, d66);
	xor (d302, d238, d255);
	and (d303, d220, d235);
	nor (d304, d223, d242);
	not (d305, d211);
	and (d306, d214, d247);
	buf (d307, d1);
	buf (d308, d138);
	not (d309, d140);
	nand (d310, d239, d243);
	nor (d311, d244, d251);
	not (d312, d100);
	buf (d313, d194);
	nor (d314, d234, d244);
	nand (d315, d234, d244);
	buf (d316, d184);
	or (d317, d212, d217);
	not (d318, d43);
	nand (d319, d210, d246);
	xor (d320, d225, d228);
	not (d321, d128);
	buf (d322, d149);
	nand (d323, d217, d252);
	xnor (d324, d219);
	and (d325, d221, d240);
	nor (d326, d235, d247);
	nand (d327, d294, d303);
	xor (d328, d273, d280);
	not (d329, d177);
	buf (d330, d225);
	not (d331, d88);
	nand (d332, d289, d326);
	buf (d333, d241);
	xnor (d334, d310, d317);
	xor (d335, d264, d274);
	not (d336, d267);
	nand (d337, d263, d307);
	xor (d338, d299, d315);
	xnor (d339, d266, d268);
	xnor (d340, d290, d306);
	not (d341, d105);
	xnor (d342, d264, d326);
	buf (d343, d2);
	xnor (d344, d298, d323);
	nand (d345, d274, d320);
	buf (d346, d169);
	xnor (d347, d296, d323);
	xor (d348, d280);
	buf (d349, d218);
	not (d350, d269);
	and (d351, d267, d304);
	and (d352, d292, d305);
	nor (d353, d264, d279);
	nand (d354, d293, d312);
	nand (d355, d272, d274);
	xnor (d356, d259, d316);
	buf (d357, d81);
	buf (d358, d260);
	nand (d359, d258, d285);
	xnor (d360, d289, d325);
	xnor (d361, d311, d323);
	or (d362, d258, d321);
	nand (d363, d265, d312);
	or (d364, d271, d278);
	nand (d365, d258, d289);
	or (d366, d268, d310);
	buf (d367, d232);
	xnor (d368, d268, d321);
	not (d369, d301);
	not (d370, d115);
	or (d371, d269, d318);
	not (d372, d188);
	xor (d373, d295, d317);
	nand (d374, d276, d301);
	or (d375, d259, d314);
	or (d376, d271, d298);
	buf (d377, d14);
	and (d378, d319, d321);
	xnor (d379, d275, d311);
	xnor (d380, d330, d374);
	not (d381, d176);
	xor (d382, d341, d348);
	or (d383, d363, d365);
	or (d384, d359, d367);
	nor (d385, d334, d350);
	xnor (d386, d354, d367);
	nor (d387, d331, d332);
	nor (d388, d332, d338);
	nand (d389, d331, d379);
	xor (d390, d365, d375);
	nor (d391, d339, d372);
	and (d392, d327, d341);
	and (d393, d332, d379);
	and (d394, d335, d361);
	xor (d395, d354, d357);
	buf (d396, d113);
	xnor (d397, d337, d371);
	xor (d398, d367, d370);
	nand (d399, d354, d379);
	not (d400, d185);
	nand (d401, d357, d372);
	or (d402, d337, d376);
	or (d403, d335, d358);
	buf (d404, d158);
	nor (d405, d331, d373);
	not (d406, d12);
	or (d407, d332, d363);
	nand (d408, d363, d365);
	xor (d409, d355);
	not (d410, d232);
	and (d411, d334, d363);
	not (d412, d42);
	or (d413, d346, d365);
	xnor (d414, d347, d358);
	nor (d415, d348, d359);
	nand (d416, d338, d368);
	or (d417, d331, d338);
	xnor (d418, d345, d352);
	xor (d419, d336, d377);
	xnor (d420, d359, d373);
	and (d421, d330, d348);
	nor (d422, d356, d377);
	xor (d423, d327, d337);
	buf (d424, d331);
	xnor (d425, d338, d350);
	xor (d426, d369, d371);
	xnor (d427, d332, d346);
	xor (d428, d360, d372);
	nand (d429, d339, d378);
	not (d430, d131);
	xor (d431, d345);
	and (d432, d329, d351);
	nand (d433, d334, d374);
	nand (d434, d370, d375);
	nand (d435, d330, d360);
	and (d436, d365, d370);
	buf (d437, d300);
	not (d438, d97);
	or (d439, d357, d376);
	nor (d440, d342, d344);
	and (d441, d328, d365);
	xnor (d442, d339, d351);
	and (d443, d354, d364);
	and (d444, d368, d370);
	nor (d445, d340, d369);
	nand (d446, d345, d371);
	nand (d447, d358, d371);
	xor (d448, d335, d337);
	buf (d449, d32);
	or (d450, d331, d353);
	not (d451, d204);
	xnor (d452, d362, d376);
	buf (d453, d346);
	not (d454, d81);
	not (d455, d27);
	xor (d456, d332, d378);
	xnor (d457, d350, d354);
	nand (d458, d351, d355);
	nand (d459, d361, d365);
	xnor (d460, d418, d458);
	and (d461, d418, d450);
	nor (d462, d406, d424);
	nand (d463, d390, d418);
	not (d464, d418);
	not (d465, d247);
	or (d466, d416, d441);
	nor (d467, d407, d418);
	or (d468, d438, d452);
	nor (d469, d411, d420);
	xnor (d470, d388, d410);
	xor (d471, d401, d421);
	not (d472, d199);
	xor (d473, d426, d431);
	xnor (d474, d415, d439);
	buf (d475, d453);
	xor (d476, d429);
	and (d477, d388, d429);
	xnor (d478, d385, d429);
	not (d479, d158);
	or (d480, d406, d422);
	xnor (d481, d395, d456);
	nor (d482, d406, d429);
	xor (d483, d382, d417);
	buf (d484, d425);
	buf (d485, d98);
	buf (d486, d96);
	not (d487, d152);
	or (d488, d429, d433);
	xnor (d489, d420, d427);
	and (d490, d422, d433);
	buf (d491, d183);
	nor (d492, d406, d420);
	or (d493, d393, d441);
	nand (d494, d407, d449);
	nor (d495, d427, d448);
	buf (d496, d185);
	nor (d497, d418, d450);
	xnor (d498, d409, d429);
	and (d499, d395, d408);
	xnor (d500, d389, d405);
	or (d501, d390, d408);
	not (d502, d254);
	buf (d503, d376);
	and (d504, d394, d414);
	and (d505, d393, d436);
	buf (d506, d324);
	or (d507, d392, d403);
	nand (d508, d433, d442);
	or (d509, d384, d441);
	and (d510, d384, d448);
	or (d511, d380, d386);
	and (d512, d409, d421);
	and (d513, d453, d457);
	xnor (d514, d426, d430);
	xnor (d515, d399, d412);
	or (d516, d389, d430);
	or (d517, d420, d440);
	xnor (d518, d399, d443);
	nor (d519, d431, d457);
	xor (d520, d401, d415);
	nand (d521, d404, d420);
	nor (d522, d432, d454);
	nor (d523, d390, d413);
	xnor (d524, d410, d439);
	buf (d525, d269);
	not (d526, d349);
	and (d527, d393, d449);
	buf (d528, d190);
	or (d529, d410, d423);
	buf (d530, d143);
	or (d531, d423, d431);
	nor (d532, d416, d419);
	not (d533, d35);
	or (d534, d468, d475);
	xnor (d535, d471, d491);
	xor (d536, d483, d508);
	or (d537, d460, d485);
	or (d538, d508, d533);
	nor (d539, d475, d495);
	and (d540, d510, d524);
	nor (d541, d477, d525);
	and (d542, d494, d523);
	xor (d543, d482, d518);
	and (d544, d482, d497);
	xnor (d545, d509, d516);
	or (d546, d487, d523);
	xor (d547, d475, d512);
	buf (d548, d398);
	xor (d549, d499, d522);
	xnor (d550, d483, d505);
	nand (d551, d476, d506);
	nand (d552, d465, d522);
	buf (d553, d460);
	not (d554, d66);
	xor (d555, d464, d482);
	or (d556, d480, d491);
	or (d557, d465, d477);
	not (d558, d276);
	or (d559, d508, d521);
	nor (d560, d481, d520);
	xnor (d561, d477, d515);
	xnor (d562, d462, d477);
	nand (d563, d464, d497);
	xor (d564, d476, d503);
	and (d565, d462);
	xnor (d566, d463, d513);
	nand (d567, d491, d509);
	nand (d568, d487, d532);
	nand (d569, d461, d503);
	xnor (d570, d484, d520);
	assign f1 = d570;
	assign f2 = d560;
	assign f3 = d556;
	assign f4 = d546;
	assign f5 = d542;
	assign f6 = d543;
	assign f7 = d535;
	assign f8 = d541;
	assign f9 = d544;
	assign f10 = d543;
endmodule
