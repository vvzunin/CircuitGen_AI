module CCGRCG144( x0, x1, x2, x3, x4, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17 );

	input x0, x1, x2, x3, x4;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314, d315, d316, d317, d318, d319, d320, d321, d322, d323, d324, d325, d326, d327, d328, d329, d330, d331, d332, d333, d334, d335, d336, d337, d338, d339, d340, d341, d342, d343, d344, d345, d346, d347, d348, d349, d350, d351, d352, d353, d354, d355, d356, d357, d358, d359, d360, d361, d362, d363, d364, d365, d366, d367, d368, d369, d370, d371, d372, d373, d374, d375, d376, d377, d378, d379, d380, d381, d382, d383, d384, d385, d386, d387, d388, d389, d390, d391, d392, d393, d394, d395, d396, d397, d398, d399, d400, d401, d402, d403, d404, d405, d406, d407, d408, d409, d410, d411, d412, d413, d414, d415, d416, d417, d418, d419, d420, d421, d422, d423, d424, d425, d426, d427, d428, d429, d430, d431, d432, d433, d434, d435, d436, d437, d438, d439, d440, d441, d442, d443, d444, d445, d446, d447, d448, d449, d450, d451, d452, d453, d454, d455, d456, d457, d458, d459, d460, d461, d462, d463, d464, d465, d466, d467, d468, d469, d470, d471, d472, d473, d474, d475, d476, d477, d478, d479, d480, d481, d482, d483, d484, d485, d486, d487, d488, d489, d490, d491, d492, d493, d494, d495, d496, d497, d498, d499, d500, d501, d502, d503, d504, d505, d506, d507, d508, d509, d510, d511, d512, d513, d514, d515, d516, d517, d518, d519, d520, d521, d522, d523, d524, d525, d526, d527, d528, d529, d530, d531, d532, d533, d534, d535, d536, d537, d538, d539, d540, d541, d542, d543, d544, d545, d546, d547, d548, d549, d550, d551, d552, d553, d554, d555, d556;

	not (d1, x0);
	nor (d2, x0, x3);
	xor (d3, x1, x2);
	buf (d4, x4);
	not (d5, x2);
	nor (d6, x1, x2);
	or (d7, x1, x4);
	and (d8, x2, x4);
	xor (d9, x0);
	buf (d10, x0);
	nor (d11, x3, x4);
	nand (d12, x2, x4);
	buf (d13, x2);
	and (d14, x1, x2);
	nand (d15, x0, x4);
	nand (d16, x3);
	nor (d17, x3);
	nand (d18, x4);
	buf (d19, x3);
	and (d20, x2, x3);
	not (d21, x4);
	and (d22, x2, x3);
	or (d23, x1, x4);
	nand (d24, x1, x4);
	xnor (d25, x0, x3);
	or (d26, x0, x1);
	buf (d27, x1);
	or (d28, x3, x4);
	not (d29, x3);
	not (d30, x1);
	nor (d31, x0, x4);
	nand (d32, x1, x2);
	xnor (d33, x2, x3);
	xnor (d34, x1, x3);
	xnor (d35, x1, x2);
	nand (d36, x3, x4);
	nor (d37, x2, x4);
	xnor (d38, x2, x3);
	nor (d39, x0, x3);
	xor (d40, x1, x3);
	nor (d41, x1, x3);
	nand (d42, x3, x4);
	xor (d43, x0, x1);
	xnor (d44, x1, x4);
	nor (d45, x2, x3);
	nand (d46, x0, x1);
	xnor (d47, x2, x4);
	and (d48, x0, x4);
	nand (d49, x2, x3);
	xnor (d50, x2);
	nor (d51, x2, x4);
	xor (d52, x1, x4);
	nor (d53, x1);
	nor (d54, d12, d38);
	and (d55, d5, d28);
	xnor (d56, d12, d23);
	buf (d57, d4);
	not (d58, d17);
	nand (d59, d41, d47);
	xnor (d60, d8, d11);
	xnor (d61, d16, d19);
	and (d62, d16, d41);
	not (d63, d1);
	not (d64, d34);
	or (d65, d31, d53);
	not (d66, d20);
	or (d67, d7, d19);
	nor (d68, d22, d30);
	not (d69, d39);
	or (d70, d8, d46);
	not (d71, d6);
	xnor (d72, d34, d38);
	xnor (d73, d35, d42);
	and (d74, d12, d34);
	nor (d75, d37, d50);
	buf (d76, d46);
	and (d77, d29, d34);
	and (d78, d48, d53);
	not (d79, d45);
	xor (d80, d17, d35);
	nand (d81, d20, d51);
	xnor (d82, d11, d50);
	buf (d83, d21);
	buf (d84, d41);
	xnor (d85, d32, d33);
	xnor (d86, d35, d53);
	xnor (d87, d40, d49);
	or (d88, d28, d37);
	and (d89, d21, d51);
	or (d90, d20, d44);
	and (d91, d25, d33);
	nand (d92, d16, d28);
	not (d93, d15);
	nand (d94, d11, d30);
	nand (d95, d1, d46);
	nor (d96, d5, d23);
	nand (d97, d26, d53);
	nor (d98, d9, d50);
	xnor (d99, d10, d33);
	nand (d100, d6, d23);
	buf (d101, d35);
	xnor (d102, d79, d98);
	and (d103, d54, d94);
	not (d104, d78);
	nor (d105, d100);
	nand (d106, d82, d101);
	nor (d107, d64, d90);
	nand (d108, d54, d99);
	or (d109, d71, d83);
	buf (d110, d72);
	and (d111, d63, d88);
	buf (d112, d56);
	nand (d113, d70, d92);
	nor (d114, d61, d62);
	and (d115, d81, d92);
	xnor (d116, d55, d61);
	not (d117, d27);
	and (d118, d64, d67);
	not (d119, d8);
	nor (d120, d57, d71);
	xor (d121, d60, d75);
	and (d122, d68, d80);
	not (d123, d93);
	nand (d124, d56, d70);
	nand (d125, d56, d74);
	and (d126, d61, d91);
	nand (d127, d64, d67);
	and (d128, d89, d99);
	and (d129, d69, d88);
	nor (d130, d65, d85);
	nor (d131, d71, d74);
	and (d132, d59, d98);
	xnor (d133, d55, d85);
	not (d134, d67);
	xnor (d135, d87, d94);
	nor (d136, d70, d92);
	not (d137, d51);
	or (d138, d67, d91);
	or (d139, d80, d91);
	buf (d140, d90);
	or (d141, d57, d77);
	xor (d142, d58, d95);
	nand (d143, d71, d73);
	xnor (d144, d65, d69);
	or (d145, d59, d86);
	nand (d146, d55, d96);
	and (d147, d75, d87);
	xor (d148, d75, d88);
	and (d149, d61, d62);
	not (d150, d63);
	not (d151, d58);
	xor (d152, d57, d70);
	xnor (d153, d96, d98);
	and (d154, d82, d87);
	xor (d155, d55, d94);
	nor (d156, d73, d81);
	not (d157, d65);
	nor (d158, d89, d91);
	and (d159, d55, d82);
	nand (d160, d66, d93);
	buf (d161, d99);
	not (d162, d79);
	xnor (d163, d63, d84);
	xnor (d164, d57, d85);
	xor (d165, d61, d99);
	or (d166, d72, d77);
	xnor (d167, d63, d76);
	not (d168, d49);
	or (d169, d56, d70);
	nor (d170, d59, d63);
	or (d171, d56, d79);
	not (d172, d35);
	or (d173, d56, d64);
	nor (d174, d58, d60);
	nor (d175, d83, d101);
	xor (d176, d72, d91);
	buf (d177, d22);
	nor (d178, d66, d92);
	and (d179, d56, d94);
	buf (d180, d60);
	or (d181, d58, d80);
	xnor (d182, d80, d81);
	not (d183, d74);
	not (d184, d16);
	nor (d185, d61, d96);
	buf (d186, d59);
	nand (d187, d59, d85);
	not (d188, d55);
	and (d189, d86, d99);
	nand (d190, d128, d164);
	and (d191, d134, d150);
	buf (d192, d85);
	or (d193, d156, d189);
	and (d194, d107, d151);
	buf (d195, d125);
	or (d196, d183, d185);
	xor (d197, d168, d179);
	nand (d198, d127, d175);
	not (d199, d80);
	xor (d200, d135, d157);
	and (d201, d138, d168);
	nand (d202, d105, d123);
	xnor (d203, d140, d148);
	nor (d204, d113, d133);
	xor (d205, d103, d140);
	not (d206, d138);
	not (d207, d57);
	or (d208, d111, d170);
	xor (d209, d146, d149);
	nor (d210, d158, d161);
	xnor (d211, d123, d169);
	and (d212, d108, d142);
	not (d213, d163);
	buf (d214, d188);
	xor (d215, d212, d213);
	xnor (d216, d210, d211);
	buf (d217, d52);
	nand (d218, d206, d214);
	and (d219, d190, d202);
	not (d220, d119);
	and (d221, d194, d210);
	xnor (d222, d200, d209);
	or (d223, d195, d214);
	buf (d224, d12);
	nor (d225, d203, d204);
	nor (d226, d202, d208);
	or (d227, d199, d206);
	xnor (d228, d206, d210);
	xnor (d229, d202);
	xor (d230, d197, d209);
	xor (d231, d193, d207);
	buf (d232, d211);
	xor (d233, d197, d203);
	nor (d234, d201, d209);
	nand (d235, d196, d197);
	and (d236, d195, d205);
	nor (d237, d197, d205);
	and (d238, d195, d205);
	xnor (d239, d191, d209);
	xnor (d240, d190, d197);
	xnor (d241, d204, d208);
	xor (d242, d206, d211);
	and (d243, d209, d211);
	xnor (d244, d196, d209);
	or (d245, d191, d202);
	nand (d246, d205, d209);
	nor (d247, d191, d206);
	nand (d248, d196, d202);
	xnor (d249, d194, d203);
	xor (d250, d196, d202);
	xnor (d251, d195, d208);
	buf (d252, d213);
	or (d253, d190, d197);
	not (d254, d151);
	or (d255, d200, d207);
	xnor (d256, d214);
	xnor (d257, d193, d198);
	xnor (d258, d194, d205);
	xor (d259, d195, d209);
	buf (d260, d3);
	not (d261, d166);
	and (d262, d197, d210);
	xnor (d263, d192, d210);
	nand (d264, d201, d214);
	nor (d265, d205);
	or (d266, d210, d211);
	and (d267, d190, d213);
	or (d268, d203, d204);
	buf (d269, d81);
	or (d270, d209, d214);
	buf (d271, d65);
	nor (d272, d198, d212);
	nand (d273, d210, d211);
	and (d274, d204, d209);
	xor (d275, d192, d213);
	not (d276, d159);
	xnor (d277, d209);
	nor (d278, d191, d205);
	or (d279, d192, d209);
	nand (d280, d196);
	xnor (d281, d206, d207);
	nand (d282, d190, d205);
	or (d283, d204, d211);
	and (d284, d195, d201);
	and (d285, d191, d200);
	xor (d286, d234, d268);
	not (d287, d167);
	xor (d288, d216, d246);
	xnor (d289, d286, d288);
	or (d290, d287, d288);
	nand (d291, d286, d288);
	or (d292, d288);
	and (d293, d288);
	not (d294, d156);
	and (d295, d287);
	buf (d296, d140);
	buf (d297, d34);
	xnor (d298, d286, d288);
	not (d299, d288);
	not (d300, d172);
	xor (d301, d286, d287);
	and (d302, d286, d287);
	not (d303, d235);
	nor (d304, d287, d288);
	buf (d305, d93);
	nor (d306, d286, d288);
	and (d307, d286, d288);
	nand (d308, d288);
	xnor (d309, d287, d288);
	and (d310, d286);
	xor (d311, d286, d288);
	and (d312, d287, d288);
	nor (d313, d286, d287);
	or (d314, d286);
	buf (d315, d265);
	not (d316, d256);
	nor (d317, d286, d287);
	xnor (d318, d287);
	nand (d319, d286, d287);
	buf (d320, d38);
	not (d321, d118);
	xor (d322, d286);
	buf (d323, d6);
	xor (d324, d287);
	or (d325, d286, d288);
	not (d326, d10);
	buf (d327, d15);
	xor (d328, d287, d288);
	and (d329, d287, d288);
	nand (d330, d287);
	xnor (d331, d286);
	nand (d332, d286, d288);
	xor (d333, d288);
	not (d334, d37);
	nor (d335, d287);
	buf (d336, d108);
	or (d337, d291, d315);
	or (d338, d318, d321);
	buf (d339, d320);
	buf (d340, d221);
	xnor (d341, d326, d328);
	not (d342, d284);
	xor (d343, d293, d321);
	buf (d344, d230);
	xor (d345, d295, d328);
	and (d346, d289, d317);
	nand (d347, d300, d335);
	and (d348, d312, d313);
	nor (d349, d314, d318);
	xnor (d350, d307, d328);
	and (d351, d302, d335);
	xnor (d352, d301, d322);
	xnor (d353, d299, d327);
	xnor (d354, d327, d333);
	buf (d355, d276);
	not (d356, d195);
	nor (d357, d298, d299);
	xor (d358, d299, d332);
	nor (d359, d316, d331);
	or (d360, d304, d306);
	or (d361, d298, d313);
	xnor (d362, d314, d334);
	xor (d363, d315, d324);
	nor (d364, d308, d323);
	nand (d365, d302, d308);
	nor (d366, d313, d335);
	not (d367, d22);
	buf (d368, d244);
	xnor (d369, d297, d310);
	nand (d370, d294, d297);
	buf (d371, d39);
	nand (d372, d290, d320);
	or (d373, d317, d329);
	buf (d374, d123);
	or (d375, d304, d322);
	and (d376, d291, d328);
	or (d377, d311, d317);
	nor (d378, d301, d336);
	and (d379, d311, d320);
	xnor (d380, d295, d299);
	nand (d381, d293, d335);
	xor (d382, d296, d298);
	buf (d383, d19);
	xor (d384, d295, d315);
	nand (d385, d311, d332);
	and (d386, d292, d312);
	and (d387, d299, d306);
	buf (d388, d200);
	xor (d389, d292, d310);
	xnor (d390, d304, d326);
	nor (d391, d316, d319);
	not (d392, d269);
	xnor (d393, d292, d335);
	xor (d394, d309, d336);
	not (d395, d199);
	xor (d396, d301, d321);
	xor (d397, d296, d307);
	xnor (d398, d311, d317);
	xor (d399, d314, d326);
	or (d400, d311, d336);
	or (d401, d322, d331);
	or (d402, d306, d331);
	xor (d403, d292, d316);
	xor (d404, d305, d312);
	xor (d405, d303, d307);
	xor (d406, d298, d331);
	not (d407, d290);
	buf (d408, d225);
	or (d409, d317, d320);
	not (d410, d245);
	buf (d411, d261);
	or (d412, d298, d311);
	and (d413, d302, d305);
	nand (d414, d295, d315);
	nor (d415, d296, d308);
	nand (d416, d296, d301);
	not (d417, d161);
	or (d418, d294, d327);
	or (d419, d292, d328);
	nand (d420, d291, d293);
	nand (d421, d302, d329);
	nor (d422, d377, d400);
	and (d423, d340, d370);
	buf (d424, d390);
	xnor (d425, d338, d387);
	xor (d426, d409, d419);
	nor (d427, d343, d401);
	and (d428, d343, d359);
	nand (d429, d368, d370);
	or (d430, d340, d357);
	buf (d431, d363);
	xnor (d432, d366, d403);
	xor (d433, d360, d383);
	nand (d434, d387, d396);
	not (d435, d81);
	not (d436, d280);
	nor (d437, d394, d414);
	not (d438, d32);
	nand (d439, d338, d390);
	xnor (d440, d395, d398);
	nor (d441, d346, d372);
	nand (d442, d346, d398);
	buf (d443, d409);
	xnor (d444, d343, d353);
	nor (d445, d359, d408);
	xor (d446, d354, d374);
	xnor (d447, d355, d356);
	or (d448, d400, d411);
	and (d449, d359, d401);
	and (d450, d390, d393);
	xor (d451, d380, d418);
	buf (d452, d141);
	nor (d453, d358, d399);
	nand (d454, d369, d405);
	or (d455, d364, d379);
	not (d456, d143);
	buf (d457, d109);
	not (d458, d36);
	or (d459, d382, d400);
	nor (d460, d368, d374);
	nand (d461, d369, d391);
	nand (d462, d395, d421);
	nand (d463, d366, d419);
	or (d464, d360, d382);
	nor (d465, d343, d355);
	xor (d466, d338, d365);
	xor (d467, d364, d385);
	buf (d468, d235);
	xor (d469, d350, d363);
	and (d470, d341, d411);
	and (d471, d401, d416);
	xnor (d472, d351, d378);
	nor (d473, d365, d369);
	nand (d474, d380, d396);
	buf (d475, d142);
	nand (d476, d359, d366);
	xor (d477, d364, d406);
	and (d478, d358, d373);
	xnor (d479, d347, d381);
	or (d480, d362, d385);
	xnor (d481, d340, d390);
	or (d482, d354, d413);
	and (d483, d363, d371);
	xnor (d484, d375, d384);
	xor (d485, d381, d390);
	and (d486, d367);
	buf (d487, d367);
	nand (d488, d353, d355);
	nand (d489, d358, d411);
	nor (d490, d407, d419);
	buf (d491, d164);
	xor (d492, d373, d401);
	nand (d493, d374, d405);
	nand (d494, d337, d353);
	nand (d495, d381, d411);
	nor (d496, d349, d396);
	xor (d497, d388, d389);
	xnor (d498, d379, d412);
	buf (d499, d120);
	nand (d500, d337, d419);
	not (d501, d275);
	and (d502, d340, d392);
	xor (d503, d375, d385);
	or (d504, d366, d371);
	nor (d505, d338, d351);
	nand (d506, d360, d368);
	not (d507, d148);
	and (d508, d342, d347);
	xnor (d509, d344, d370);
	xor (d510, d339, d366);
	or (d511, d353, d411);
	and (d512, d366, d396);
	buf (d513, d18);
	nand (d514, d390, d410);
	xor (d515, d398, d418);
	xor (d516, d379, d391);
	buf (d517, d416);
	xor (d518, d397, d416);
	buf (d519, d351);
	xnor (d520, d439, d453);
	and (d521, d473, d480);
	or (d522, d431, d435);
	not (d523, d126);
	or (d524, d491, d507);
	not (d525, d390);
	and (d526, d512, d514);
	and (d527, d468, d516);
	buf (d528, d397);
	and (d529, d448, d495);
	nor (d530, d449, d482);
	not (d531, d500);
	not (d532, d399);
	nand (d533, d434, d514);
	or (d534, d466, d477);
	not (d535, d24);
	xnor (d536, d512, d515);
	buf (d537, d294);
	nor (d538, d440, d486);
	or (d539, d450, d500);
	not (d540, d393);
	buf (d541, d435);
	and (d542, d465, d474);
	nor (d543, d459, d487);
	and (d544, d481, d487);
	xnor (d545, d458, d460);
	nor (d546, d507, d512);
	nand (d547, d441, d498);
	xor (d548, d477, d485);
	not (d549, d219);
	nor (d550, d439, d505);
	not (d551, d43);
	xnor (d552, d438, d491);
	xnor (d553, d493, d515);
	nand (d554, d466, d493);
	or (d555, d462, d491);
	and (d556, d437, d453);
	assign f1 = d549;
	assign f2 = d549;
	assign f3 = d545;
	assign f4 = d525;
	assign f5 = d524;
	assign f6 = d530;
	assign f7 = d536;
	assign f8 = d551;
	assign f9 = d541;
	assign f10 = d543;
	assign f11 = d543;
	assign f12 = d550;
	assign f13 = d530;
	assign f14 = d551;
	assign f15 = d533;
	assign f16 = d530;
	assign f17 = d529;
endmodule
