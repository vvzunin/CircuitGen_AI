module CCGRCG75( x0, x1, x2, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17, f18, f19, f20 );

	input x0, x1, x2;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17, f18, f19, f20;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314, d315, d316, d317, d318, d319, d320, d321, d322, d323, d324, d325, d326, d327, d328, d329, d330, d331, d332, d333, d334, d335, d336, d337, d338, d339, d340, d341, d342, d343, d344, d345, d346, d347, d348, d349, d350, d351, d352, d353, d354, d355, d356, d357, d358, d359, d360, d361, d362, d363, d364, d365, d366, d367, d368, d369, d370, d371, d372, d373, d374, d375, d376, d377, d378, d379, d380, d381, d382, d383, d384, d385, d386, d387, d388, d389, d390, d391, d392, d393, d394, d395, d396, d397, d398, d399, d400, d401, d402, d403, d404, d405, d406, d407, d408, d409, d410, d411, d412, d413, d414, d415, d416, d417, d418, d419, d420, d421, d422, d423, d424, d425, d426, d427, d428, d429, d430;

	xor (d1, x1);
	not (d2, x0);
	nand (d3, x0, x2);
	nor (d4, x0, x1);
	or (d5, x2);
	nand (d6, x0);
	not (d7, x2);
	and (d8, x0, x1);
	or (d9, d1, d3);
	buf (d10, x1);
	buf (d11, x0);
	not (d12, d6);
	xnor (d13, d4, d5);
	xnor (d14, d2, d7);
	nand (d15, d6, d8);
	nand (d16, d2, d6);
	nor (d17, d4, d5);
	xnor (d18, d8);
	or (d19, d4, d6);
	xnor (d20, d2, d4);
	nand (d21, d5);
	or (d22, d5, d6);
	buf (d23, d2);
	not (d24, d1);
	buf (d25, d6);
	xnor (d26, d7, d8);
	buf (d27, d5);
	xnor (d28, d1, d8);
	and (d29, d6, d7);
	or (d30, d6, d7);
	nor (d31, d3, d7);
	and (d32, d1, d3);
	and (d33, d7, d8);
	nand (d34, d1, d2);
	nand (d35, d1, d6);
	and (d36, d1, d4);
	or (d37, d4, d6);
	buf (d38, d1);
	and (d39, d1, d7);
	xor (d40, d4, d8);
	and (d41, d1, d7);
	nor (d42, d7);
	or (d43, d7, d8);
	or (d44, d4, d8);
	xor (d45, d5, d7);
	nand (d46, d4, d7);
	xor (d47, d4, d6);
	buf (d48, d8);
	nand (d49, d2, d8);
	and (d50, d3, d8);
	xor (d51, d2, d6);
	xor (d52, d3, d8);
	and (d53, d4);
	xnor (d54, d1, d7);
	nor (d55, d2, d6);
	or (d56, d2, d8);
	nor (d57, d7, d8);
	xnor (d58, d4, d7);
	and (d59, d1, d2);
	buf (d60, d4);
	and (d61, d1, d6);
	xor (d62, d1);
	nand (d63, d2, d3);
	or (d64, d3, d6);
	buf (d65, d7);
	nand (d66, d1, d5);
	xor (d67, d7, d8);
	xnor (d68, d4, d6);
	nand (d69, d2, d8);
	not (d70, d65);
	nor (d71, d19, d50);
	nand (d72, d19, d41);
	nand (d73, d30, d59);
	not (d74, d69);
	nor (d75, d28, d61);
	buf (d76, d25);
	xnor (d77, d24, d49);
	not (d78, d26);
	xor (d79, d12, d40);
	or (d80, d22, d65);
	nor (d81, d61, d63);
	xnor (d82, d54, d57);
	and (d83, d54, d55);
	nor (d84, d17, d39);
	nor (d85, d34, d52);
	or (d86, d57, d60);
	xor (d87, d28, d51);
	nand (d88, d19, d31);
	or (d89, d45, d55);
	xor (d90, d39, d63);
	nor (d91, d20, d55);
	or (d92, d42, d61);
	or (d93, d48, d69);
	nand (d94, d28, d50);
	xor (d95, d44, d67);
	nand (d96, d38, d64);
	not (d97, d34);
	xnor (d98, d23, d53);
	xor (d99, d13, d53);
	nand (d100, d21, d42);
	not (d101, d24);
	buf (d102, d33);
	nor (d103, d60, d69);
	nor (d104, d29, d35);
	xor (d105, d35, d54);
	xor (d106, d29, d65);
	xor (d107, d14, d16);
	xnor (d108, d30, d34);
	xor (d109, d21, d55);
	xor (d110, d62, d63);
	not (d111, d43);
	not (d112, d27);
	xnor (d113, d15, d63);
	and (d114, d33, d67);
	nand (d115, d10, d65);
	nand (d116, d21, d27);
	xnor (d117, d16, d18);
	and (d118, d43, d44);
	not (d119, d30);
	and (d120, d56, d57);
	xnor (d121, d44, d64);
	or (d122, d23, d64);
	and (d123, d29, d34);
	xor (d124, d25, d32);
	not (d125, d9);
	not (d126, d38);
	buf (d127, d39);
	nand (d128, d24, d56);
	or (d129, d31, d66);
	buf (d130, d38);
	nand (d131, d12, d61);
	nor (d132, d39, d41);
	xnor (d133, d33, d66);
	nand (d134, d14, d17);
	nor (d135, d32, d63);
	and (d136, d61, d69);
	or (d137, d17, d44);
	and (d138, d49, d58);
	xor (d139, d48, d56);
	nand (d140, d43, d47);
	nand (d141, d13, d20);
	not (d142, d56);
	xnor (d143, d13, d63);
	or (d144, d13, d60);
	or (d145, d32, d68);
	buf (d146, d13);
	not (d147, d62);
	nand (d148, d28, d44);
	or (d149, d24, d65);
	xor (d150, d58, d68);
	or (d151, d11, d27);
	xor (d152, d36, d48);
	or (d153, d69);
	or (d154, d12, d21);
	or (d155, d48, d51);
	xor (d156, d34, d57);
	buf (d157, d28);
	xnor (d158, d89, d111);
	nor (d159, d72, d137);
	xnor (d160, d151, d153);
	xnor (d161, d160);
	not (d162, d146);
	xor (d163, d158);
	or (d164, d158, d159);
	buf (d165, d54);
	buf (d166, d3);
	and (d167, d159, d160);
	nor (d168, d159, d160);
	nand (d169, d162, d167);
	buf (d170, d151);
	or (d171, d163, d167);
	xor (d172, d161, d163);
	nand (d173, d162, d168);
	not (d174, d156);
	nand (d175, d165, d167);
	and (d176, d165, d168);
	not (d177, d11);
	xnor (d178, d162, d164);
	or (d179, d161, d163);
	xnor (d180, d162, d163);
	nor (d181, d164);
	buf (d182, d30);
	xnor (d183, d162, d168);
	or (d184, d162, d168);
	buf (d185, d98);
	and (d186, d166, d167);
	nand (d187, d164, d168);
	xor (d188, d162, d165);
	nor (d189, d165, d168);
	and (d190, d161, d163);
	nand (d191, d162);
	xor (d192, d162, d165);
	nor (d193, d162, d168);
	buf (d194, d83);
	buf (d195, d155);
	nand (d196, d164);
	xor (d197, d161, d162);
	xor (d198, d161, d168);
	xor (d199, d163, d164);
	or (d200, d165, d168);
	nand (d201, d166, d168);
	nor (d202, d162);
	xor (d203, d164, d166);
	and (d204, d162, d165);
	buf (d205, d152);
	buf (d206, d51);
	nand (d207, d162, d165);
	and (d208, d164, d167);
	xor (d209, d165, d168);
	nor (d210, d163, d164);
	buf (d211, d47);
	or (d212, d163, d166);
	nor (d213, d162, d167);
	xor (d214, d166, d168);
	or (d215, d179, d181);
	nand (d216, d184, d199);
	nor (d217, d177, d180);
	and (d218, d176, d184);
	xnor (d219, d201, d212);
	xor (d220, d187, d198);
	or (d221, d185, d210);
	and (d222, d200, d204);
	or (d223, d200, d202);
	not (d224, d210);
	xor (d225, d193, d201);
	xor (d226, d176, d184);
	buf (d227, d208);
	xor (d228, d184, d208);
	xnor (d229, d179, d196);
	xor (d230, d169, d175);
	xor (d231, d199);
	or (d232, d188, d212);
	or (d233, d193, d208);
	nor (d234, d170, d192);
	nand (d235, d177, d209);
	nor (d236, d207, d212);
	nand (d237, d172, d186);
	buf (d238, d195);
	xor (d239, d178, d206);
	buf (d240, d62);
	buf (d241, d88);
	or (d242, d175, d191);
	nand (d243, d188, d194);
	xor (d244, d185, d214);
	xnor (d245, d196, d210);
	nor (d246, d189, d196);
	buf (d247, d211);
	buf (d248, d57);
	xnor (d249, d171, d211);
	buf (d250, d76);
	xnor (d251, d192, d200);
	xnor (d252, d197, d208);
	or (d253, d180, d195);
	nor (d254, d207, d213);
	buf (d255, d36);
	xnor (d256, d198, d200);
	xor (d257, d170, d206);
	and (d258, d206, d214);
	and (d259, d173, d190);
	nand (d260, d210);
	nand (d261, d176, d178);
	buf (d262, d67);
	nand (d263, d169, d208);
	buf (d264, d90);
	xor (d265, d214);
	and (d266, d171, d189);
	nand (d267, d170, d187);
	not (d268, d109);
	nand (d269, d182, d205);
	nor (d270, d204, d209);
	nand (d271, d212, d214);
	not (d272, d138);
	not (d273, d61);
	xor (d274, d195, d200);
	or (d275, d189, d192);
	xor (d276, d195, d214);
	or (d277, d170, d210);
	or (d278, d208, d209);
	nand (d279, d206, d207);
	xor (d280, d179, d207);
	buf (d281, d92);
	or (d282, d184, d207);
	xor (d283, d192, d194);
	and (d284, d171, d185);
	nor (d285, d170, d193);
	buf (d286, d160);
	nand (d287, d169, d213);
	and (d288, d172, d196);
	nor (d289, d199, d209);
	xnor (d290, d194, d196);
	and (d291, d242, d281);
	buf (d292, d154);
	and (d293, d238, d243);
	nand (d294, d219, d258);
	and (d295, d271, d289);
	buf (d296, d133);
	and (d297, d226, d245);
	not (d298, d132);
	buf (d299, d107);
	nand (d300, d221, d226);
	xnor (d301, d273);
	or (d302, d216, d231);
	nor (d303, d223, d234);
	buf (d304, d102);
	not (d305, d126);
	nand (d306, d219, d237);
	xor (d307, d256, d268);
	buf (d308, d241);
	xnor (d309, d260, d265);
	or (d310, d266, d273);
	nor (d311, d250, d278);
	not (d312, d18);
	xor (d313, d261, d262);
	xnor (d314, d262, d264);
	xnor (d315, d224, d275);
	nand (d316, d252, d273);
	buf (d317, d153);
	xor (d318, d230, d248);
	nand (d319, d234, d245);
	buf (d320, d198);
	and (d321, d222, d223);
	not (d322, d242);
	xnor (d323, d215, d248);
	or (d324, d275, d277);
	buf (d325, d260);
	and (d326, d219, d253);
	nand (d327, d221, d255);
	not (d328, d182);
	xor (d329, d250, d259);
	and (d330, d225, d241);
	nand (d331, d255, d275);
	nor (d332, d232, d288);
	and (d333, d236, d287);
	not (d334, d119);
	nand (d335, d219, d226);
	not (d336, d287);
	nor (d337, d221, d244);
	or (d338, d252, d254);
	not (d339, d89);
	buf (d340, d115);
	buf (d341, d137);
	xor (d342, d326, d328);
	xor (d343, d303, d315);
	xnor (d344, d334, d337);
	not (d345, d301);
	not (d346, d92);
	xor (d347, d295, d330);
	nand (d348, d305, d321);
	nor (d349, d300, d320);
	not (d350, d159);
	xor (d351, d300, d315);
	or (d352, d303, d325);
	nor (d353, d295, d300);
	not (d354, d58);
	buf (d355, d276);
	and (d356, d297, d329);
	nand (d357, d300, d313);
	nand (d358, d291, d313);
	nand (d359, d305, d316);
	buf (d360, d277);
	buf (d361, d269);
	nor (d362, d294, d327);
	buf (d363, d143);
	not (d364, d349);
	xor (d365, d361);
	nand (d366, d346, d352);
	nand (d367, d349);
	nor (d368, d353, d357);
	and (d369, d342, d349);
	not (d370, d319);
	not (d371, d53);
	nor (d372, d343, d351);
	xnor (d373, d341, d351);
	buf (d374, d173);
	nand (d375, d343, d349);
	nor (d376, d344, d348);
	or (d377, d345, d352);
	and (d378, d354, d358);
	xnor (d379, d355, d360);
	or (d380, d352, d355);
	nor (d381, d355, d356);
	xnor (d382, d349, d352);
	buf (d383, d148);
	xnor (d384, d348, d349);
	and (d385, d344, d357);
	xor (d386, d343, d355);
	nor (d387, d354, d361);
	nor (d388, d346, d355);
	xnor (d389, d343);
	and (d390, d359, d360);
	nor (d391, d353, d362);
	or (d392, d354, d358);
	xor (d393, d341, d362);
	and (d394, d353, d354);
	nand (d395, d360, d361);
	or (d396, d346, d359);
	nand (d397, d350, d353);
	nor (d398, d344, d359);
	nor (d399, d360, d361);
	xnor (d400, d355, d357);
	nand (d401, d353);
	nand (d402, d352, d357);
	not (d403, d29);
	xor (d404, d342, d350);
	nand (d405, d357, d362);
	xnor (d406, d352, d362);
	and (d407, d348, d357);
	or (d408, d347);
	and (d409, d340, d341);
	or (d410, d345, d360);
	nor (d411, d348, d358);
	nand (d412, d347, d356);
	or (d413, d348, d359);
	buf (d414, d124);
	xnor (d415, d340, d353);
	not (d416, d270);
	nand (d417, d351, d361);
	nand (d418, d354, d359);
	and (d419, d348, d358);
	nor (d420, d347, d353);
	xnor (d421, d350, d351);
	nor (d422, d340, d361);
	and (d423, d342, d350);
	and (d424, d341, d344);
	nand (d425, d352, d358);
	nand (d426, d345, d350);
	or (d427, d342, d344);
	or (d428, d341, d355);
	xor (d429, d353, d356);
	buf (d430, d329);
	assign f1 = d412;
	assign f2 = d404;
	assign f3 = d408;
	assign f4 = d423;
	assign f5 = d414;
	assign f6 = d412;
	assign f7 = d397;
	assign f8 = d394;
	assign f9 = d397;
	assign f10 = d421;
	assign f11 = d422;
	assign f12 = d377;
	assign f13 = d424;
	assign f14 = d371;
	assign f15 = d395;
	assign f16 = d412;
	assign f17 = d383;
	assign f18 = d384;
	assign f19 = d375;
	assign f20 = d368;
endmodule
