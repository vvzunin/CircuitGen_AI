module CCGRCG137( x0, x1, x2, x3, x4, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13 );

	input x0, x1, x2, x3, x4;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314, d315, d316, d317, d318, d319, d320, d321, d322, d323, d324, d325, d326, d327, d328, d329, d330, d331, d332, d333, d334, d335, d336, d337, d338, d339, d340, d341, d342, d343, d344, d345, d346, d347, d348, d349, d350, d351, d352, d353, d354, d355, d356, d357, d358, d359, d360, d361, d362, d363, d364, d365, d366, d367, d368, d369, d370, d371, d372, d373, d374, d375, d376, d377, d378, d379, d380, d381, d382, d383, d384, d385, d386, d387, d388, d389, d390, d391, d392, d393, d394, d395, d396, d397, d398, d399, d400, d401, d402, d403, d404, d405, d406, d407, d408, d409, d410, d411, d412, d413, d414, d415, d416, d417, d418, d419, d420, d421, d422, d423, d424, d425, d426, d427, d428, d429, d430, d431, d432, d433, d434, d435, d436, d437, d438, d439, d440, d441, d442, d443, d444, d445, d446, d447, d448, d449, d450, d451, d452, d453, d454;

	xor (d1, x4);
	nor (d2, x0, x4);
	xnor (d3, x4);
	not (d4, x4);
	or (d5, x0, x4);
	and (d6, x1, x4);
	and (d7, x4);
	buf (d8, x0);
	xor (d9, x0, x1);
	or (d10, x1, x3);
	buf (d11, x1);
	not (d12, x3);
	or (d13, x3, x4);
	or (d14, x1, x3);
	nand (d15, x1);
	xor (d16, x3, x4);
	and (d17, x1, x4);
	and (d18, x0, x4);
	and (d19, x3, x4);
	xor (d20, x1, x4);
	xnor (d21, x0, x2);
	nand (d22, x1, x4);
	xor (d23, x1, x3);
	xnor (d24, x2, x3);
	nor (d25, x2, x4);
	and (d26, x2, x3);
	nand (d27, x0, x4);
	and (d28, x2, x3);
	xnor (d29, x3, x4);
	xor (d30, x2, x4);
	buf (d31, x3);
	and (d32, x0, x1);
	xnor (d33, x0);
	not (d34, x2);
	buf (d35, x4);
	or (d36, x0, x1);
	nor (d37, x1);
	nor (d38, x3, x4);
	and (d39, x0, x1);
	or (d40, d24, d27);
	or (d41, d16, d22);
	xnor (d42, d22);
	nand (d43, d25, d31);
	buf (d44, d36);
	or (d45, d15, d30);
	nor (d46, d18, d19);
	nand (d47, d8, d25);
	xor (d48, d5, d37);
	nand (d49, d37, d39);
	not (d50, d26);
	buf (d51, x2);
	xor (d52, d4);
	nor (d53, d21, d24);
	not (d54, d16);
	nand (d55, d27, d37);
	xnor (d56, d9, d24);
	xor (d57, d24, d36);
	not (d58, d9);
	xnor (d59, d9, d21);
	xor (d60, d25, d28);
	xor (d61, d35, d38);
	not (d62, d8);
	xor (d63, d8, d27);
	xor (d64, d19, d20);
	or (d65, d18, d27);
	nor (d66, d15, d18);
	buf (d67, d30);
	nand (d68, d26, d36);
	xnor (d69, d15, d34);
	or (d70, d15, d36);
	xor (d71, d32, d34);
	and (d72, d10, d26);
	xor (d73, d8, d12);
	buf (d74, d23);
	and (d75, d12, d27);
	buf (d76, d7);
	nor (d77, d5, d32);
	xnor (d78, d7, d8);
	xor (d79, d19, d30);
	nor (d80, d11, d32);
	not (d81, d5);
	xnor (d82, d10, d27);
	nand (d83, d21, d28);
	xnor (d84, d15, d20);
	or (d85, d4, d13);
	not (d86, d15);
	nor (d87, d16, d39);
	nor (d88, d21, d34);
	buf (d89, d2);
	nor (d90, d3, d16);
	or (d91, d31, d36);
	or (d92, d10, d36);
	nand (d93, d21, d34);
	nand (d94, d52, d89);
	xor (d95, d46, d62);
	xor (d96, d50, d73);
	xor (d97, d65, d71);
	nor (d98, d50, d89);
	nand (d99, d49, d93);
	xnor (d100, d61, d79);
	or (d101, d52, d56);
	buf (d102, d48);
	nor (d103, d79, d83);
	nand (d104, d59, d74);
	buf (d105, d73);
	nand (d106, d95, d96);
	and (d107, d100, d103);
	and (d108, d96, d98);
	not (d109, d20);
	and (d110, d95, d101);
	buf (d111, d53);
	xnor (d112, d101, d102);
	xor (d113, d102);
	not (d114, d52);
	xor (d115, d100, d102);
	and (d116, d100, d101);
	and (d117, d95, d97);
	xor (d118, d98, d102);
	not (d119, d42);
	not (d120, d101);
	nand (d121, d101, d103);
	xnor (d122, d95, d102);
	buf (d123, d101);
	or (d124, d98, d100);
	nor (d125, d97, d101);
	xor (d126, d94, d98);
	xor (d127, d97, d99);
	or (d128, d103, d104);
	not (d129, d13);
	xnor (d130, d95, d98);
	nor (d131, d95, d97);
	buf (d132, d20);
	and (d133, d97, d102);
	xnor (d134, d98, d99);
	buf (d135, d93);
	not (d136, d32);
	xor (d137, d99, d104);
	nor (d138, d100, d101);
	xor (d139, d96, d104);
	or (d140, d94, d97);
	or (d141, d94, d104);
	xnor (d142, d95, d100);
	xnor (d143, d95, d103);
	buf (d144, d81);
	xnor (d145, d98, d101);
	xor (d146, d99, d103);
	xor (d147, d97, d101);
	nand (d148, d95);
	nor (d149, d95, d101);
	and (d150, d96, d97);
	xor (d151, d100, d104);
	nand (d152, d96, d98);
	nor (d153, d97, d99);
	xnor (d154, d94, d97);
	xor (d155, d102, d104);
	nand (d156, d101, d103);
	xor (d157, d97, d99);
	xnor (d158, d97, d98);
	nor (d159, d96, d101);
	xnor (d160, d96, d98);
	nor (d161, d102, d104);
	nand (d162, d98, d100);
	nor (d163, d94, d98);
	buf (d164, d62);
	xnor (d165, d96, d100);
	nand (d166, d96, d97);
	and (d167, d123, d134);
	nand (d168, d107, d147);
	xor (d169, d147, d159);
	xor (d170, d130, d145);
	xnor (d171, d116, d139);
	buf (d172, d156);
	nand (d173, d114, d147);
	not (d174, d145);
	buf (d175, d59);
	nand (d176, d125, d135);
	xor (d177, d112, d147);
	xor (d178, d115, d150);
	nand (d179, d109, d153);
	or (d180, d120, d162);
	and (d181, d115, d162);
	nand (d182, d112, d113);
	xnor (d183, d134, d139);
	buf (d184, d38);
	not (d185, d60);
	buf (d186, d154);
	xnor (d187, d109, d111);
	nor (d188, d141, d143);
	xor (d189, d107, d157);
	and (d190, d123, d155);
	and (d191, d131, d143);
	nor (d192, d110, d157);
	or (d193, d110, d138);
	not (d194, d69);
	not (d195, d85);
	nand (d196, d126, d127);
	xor (d197, d115, d159);
	xnor (d198, d111, d165);
	nor (d199, d138, d150);
	and (d200, d107, d162);
	buf (d201, d151);
	nand (d202, d115, d143);
	xor (d203, d109, d146);
	nand (d204, d121, d155);
	nand (d205, d107, d149);
	nor (d206, d133, d140);
	or (d207, d127, d160);
	xor (d208, d116, d133);
	or (d209, d116, d133);
	and (d210, d117, d159);
	and (d211, d151, d157);
	xor (d212, d109, d131);
	xor (d213, d115, d155);
	not (d214, d136);
	not (d215, d14);
	nand (d216, d110, d130);
	nor (d217, d112, d127);
	and (d218, d114, d164);
	xnor (d219, d142, d152);
	nand (d220, d132, d158);
	or (d221, d127, d145);
	nor (d222, d106, d107);
	and (d223, d107, d148);
	and (d224, d135, d165);
	nand (d225, d125, d163);
	buf (d226, d16);
	buf (d227, d163);
	buf (d228, d149);
	and (d229, d108, d159);
	nor (d230, d123, d148);
	or (d231, d106, d134);
	xnor (d232, d113, d144);
	and (d233, d113, d124);
	buf (d234, d4);
	nor (d235, d127, d152);
	nand (d236, d148, d164);
	xor (d237, d117, d164);
	or (d238, d126, d161);
	nor (d239, d111, d136);
	xnor (d240, d115, d153);
	not (d241, d44);
	xnor (d242, d121, d164);
	xnor (d243, d119, d125);
	or (d244, d127, d141);
	buf (d245, d152);
	xor (d246, d136, d140);
	and (d247, d135, d138);
	nand (d248, d130, d135);
	xnor (d249, d198, d229);
	not (d250, d152);
	or (d251, d177, d208);
	nand (d252, d175, d244);
	xor (d253, d222, d230);
	buf (d254, d32);
	or (d255, d214, d239);
	and (d256, d215, d248);
	and (d257, d203, d233);
	xor (d258, d206, d247);
	or (d259, d167, d217);
	xor (d260, d191, d232);
	nand (d261, d185, d235);
	nand (d262, d176, d212);
	xnor (d263, d174, d177);
	not (d264, d123);
	not (d265, d25);
	and (d266, d220, d243);
	and (d267, d178, d245);
	xnor (d268, d176, d194);
	or (d269, d217, d224);
	xnor (d270, d181, d226);
	xnor (d271, d172, d226);
	or (d272, d192, d232);
	nand (d273, d256, d267);
	or (d274, d252, d256);
	xnor (d275, d249, d269);
	xor (d276, d262, d269);
	and (d277, d256, d266);
	and (d278, d261, d272);
	or (d279, d258, d261);
	xnor (d280, d260, d263);
	buf (d281, d133);
	buf (d282, d164);
	and (d283, d258, d270);
	buf (d284, d148);
	not (d285, d140);
	xor (d286, d270, d271);
	nor (d287, d254, d268);
	not (d288, d240);
	xnor (d289, d259, d261);
	xnor (d290, d258, d260);
	xor (d291, d254, d258);
	and (d292, d263, d264);
	nand (d293, d264, d265);
	nand (d294, d262, d267);
	and (d295, d249, d258);
	xnor (d296, d259, d268);
	nand (d297, d269, d270);
	not (d298, d114);
	nand (d299, d250, d269);
	nand (d300, d253, d269);
	and (d301, d252, d268);
	xnor (d302, d258, d272);
	xnor (d303, d268, d269);
	or (d304, d258, d260);
	buf (d305, d71);
	or (d306, d256, d268);
	and (d307, d263, d264);
	not (d308, d204);
	buf (d309, d79);
	xor (d310, d255, d257);
	nand (d311, d255, d261);
	xnor (d312, d255, d262);
	or (d313, d265, d270);
	and (d314, d251);
	xor (d315, d258, d259);
	and (d316, d249, d252);
	or (d317, d249, d256);
	nand (d318, d260, d266);
	nand (d319, d259, d266);
	buf (d320, d244);
	and (d321, d255, d257);
	or (d322, d249, d263);
	xnor (d323, d255, d269);
	xnor (d324, d262, d267);
	not (d325, d172);
	or (d326, d259, d261);
	or (d327, d260, d263);
	nand (d328, d251, d263);
	nor (d329, d256, d261);
	xnor (d330, d250, d263);
	or (d331, d255, d258);
	and (d332, d315, d330);
	or (d333, d299, d315);
	xor (d334, d287, d316);
	nor (d335, d278, d313);
	and (d336, d305, d324);
	and (d337, d282, d302);
	xnor (d338, d331);
	and (d339, d275, d321);
	nand (d340, d309, d316);
	xnor (d341, d278, d312);
	xnor (d342, d287, d322);
	not (d343, d174);
	buf (d344, d88);
	xor (d345, d279, d284);
	xor (d346, d296, d303);
	not (d347, d153);
	buf (d348, d12);
	nor (d349, d282, d322);
	xor (d350, d306, d329);
	nand (d351, d283, d330);
	or (d352, d287, d314);
	not (d353, d100);
	and (d354, d283, d284);
	nand (d355, d323, d329);
	or (d356, d289, d326);
	nand (d357, d280, d296);
	buf (d358, d171);
	nor (d359, d277, d285);
	xor (d360, d306, d328);
	or (d361, d287, d315);
	nand (d362, d334, d344);
	nor (d363, d340, d341);
	buf (d364, d275);
	or (d365, d347, d348);
	and (d366, d334, d348);
	buf (d367, d91);
	nor (d368, d349, d360);
	xor (d369, d355, d357);
	nand (d370, d334, d346);
	xnor (d371, d338, d353);
	xnor (d372, d337, d359);
	and (d373, d338, d345);
	not (d374, d305);
	nand (d375, d337, d354);
	nand (d376, d339, d357);
	xnor (d377, d344, d353);
	xor (d378, d347, d356);
	xnor (d379, d333, d344);
	nor (d380, d349, d359);
	xor (d381, d348, d357);
	nor (d382, d332, d343);
	or (d383, d335, d353);
	xor (d384, d334, d343);
	xor (d385, d335, d341);
	buf (d386, d102);
	xor (d387, d347, d350);
	or (d388, d335, d347);
	xor (d389, d332, d343);
	xnor (d390, d333, d354);
	or (d391, d341, d343);
	or (d392, d338, d344);
	nor (d393, d355, d357);
	not (d394, d337);
	buf (d395, d125);
	xnor (d396, d376, d390);
	and (d397, d365, d386);
	buf (d398, d331);
	not (d399, d287);
	nor (d400, d379);
	and (d401, d375, d393);
	xor (d402, d394, d395);
	nor (d403, d372, d376);
	nor (d404, d366, d384);
	nand (d405, d383, d393);
	nor (d406, d370, d385);
	buf (d407, d251);
	xor (d408, d380, d389);
	xor (d409, d372, d375);
	nand (d410, d375, d390);
	and (d411, d367, d381);
	not (d412, d281);
	nand (d413, d387, d394);
	buf (d414, d216);
	nand (d415, d383, d395);
	nor (d416, d366, d394);
	nand (d417, d382, d384);
	nand (d418, d366, d378);
	and (d419, d363, d380);
	or (d420, d365, d387);
	nor (d421, d368, d383);
	or (d422, d367, d380);
	and (d423, d370, d374);
	buf (d424, d301);
	nand (d425, d366, d388);
	and (d426, d364, d394);
	xnor (d427, d366, d378);
	and (d428, d364, d371);
	or (d429, d369, d374);
	nand (d430, d368, d389);
	xnor (d431, d377, d382);
	nor (d432, d367, d394);
	or (d433, d374, d377);
	nor (d434, d376, d384);
	buf (d435, d22);
	not (d436, d157);
	and (d437, d365, d375);
	nor (d438, d367, d368);
	xnor (d439, d370, d391);
	xnor (d440, d389, d395);
	or (d441, d373, d389);
	xnor (d442, d380, d382);
	xor (d443, d371, d381);
	nand (d444, d367, d383);
	or (d445, d376, d387);
	nand (d446, d366, d377);
	xnor (d447, d363, d375);
	not (d448, d368);
	nor (d449, d369, d378);
	xor (d450, d368, d384);
	nand (d451, d375, d383);
	nor (d452, d362, d369);
	or (d453, d362, d393);
	xnor (d454, d372, d380);
	assign f1 = d402;
	assign f2 = d428;
	assign f3 = d397;
	assign f4 = d438;
	assign f5 = d449;
	assign f6 = d447;
	assign f7 = d443;
	assign f8 = d417;
	assign f9 = d405;
	assign f10 = d427;
	assign f11 = d405;
	assign f12 = d450;
	assign f13 = d411;
endmodule
