module CCGRCG50( x0, x1, x2, f1, f2, f3, f4, f5, f6, f7, f8 );

	input x0, x1, x2;
	output f1, f2, f3, f4, f5, f6, f7, f8;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314, d315, d316, d317, d318, d319, d320, d321, d322, d323, d324, d325, d326, d327, d328, d329, d330, d331, d332, d333, d334, d335, d336, d337, d338, d339, d340, d341, d342, d343, d344, d345, d346, d347, d348, d349, d350, d351, d352, d353, d354, d355;

	and (d1, x0, x1);
	not (d2, x1);
	xnor (d3, x0, x2);
	and (d4, x0, x2);
	nand (d5, x1, x2);
	nor (d6, x0, x2);
	or (d7, x1, x2);
	buf (d8, x1);
	and (d9, x0, x1);
	and (d10, x1, x2);
	or (d11, x0, x2);
	or (d12, x0, x2);
	buf (d13, x0);
	not (d14, x0);
	xnor (d15, d1, d14);
	and (d16, d1, d12);
	nor (d17, d3, d8);
	and (d18, d6, d7);
	or (d19, d2, d11);
	xnor (d20, d1, d9);
	xor (d21, d12, d14);
	and (d22, d6, d9);
	and (d23, d11, d12);
	and (d24, d19, d21);
	nand (d25, d22);
	xnor (d26, d15, d23);
	buf (d27, d12);
	and (d28, d16, d17);
	not (d29, d21);
	buf (d30, d5);
	nand (d31, d16, d18);
	and (d32, d17, d22);
	nor (d33, d15, d21);
	nor (d34, d18, d19);
	buf (d35, d11);
	not (d36, d6);
	or (d37, d19, d21);
	not (d38, d15);
	not (d39, d2);
	xnor (d40, d19, d23);
	nor (d41, d18, d19);
	nand (d42, d19, d21);
	xnor (d43, d16, d20);
	xor (d44, d16, d22);
	xor (d45, d18, d21);
	nand (d46, d16);
	or (d47, d17, d19);
	buf (d48, d7);
	nor (d49, d17, d18);
	xnor (d50, d15, d16);
	xnor (d51, d18, d19);
	xor (d52, d16, d21);
	xnor (d53, d20, d22);
	not (d54, d20);
	nand (d55, d15, d16);
	xor (d56, d18, d22);
	buf (d57, d15);
	and (d58, d15, d17);
	nand (d59, d15, d21);
	xor (d60, d22, d23);
	nor (d61, d16, d22);
	nor (d62, d20, d21);
	xnor (d63, d17, d22);
	nor (d64, d17, d21);
	xor (d65, d57, d60);
	and (d66, d46, d55);
	and (d67, d30, d43);
	xor (d68, d32, d45);
	xnor (d69, d31, d61);
	buf (d70, d26);
	xor (d71, d39, d60);
	or (d72, d38, d41);
	buf (d73, d46);
	buf (d74, d24);
	xnor (d75, d36, d46);
	xor (d76, d26, d48);
	and (d77, d42, d53);
	nor (d78, d40, d56);
	or (d79, d27, d29);
	or (d80, d32, d40);
	nor (d81, d28, d55);
	and (d82, d36, d39);
	and (d83, d44, d60);
	nor (d84, d72, d75);
	xnor (d85, d74, d80);
	nor (d86, d76, d81);
	nor (d87, d80, d82);
	not (d88, d67);
	or (d89, d82, d83);
	buf (d90, d34);
	nand (d91, d65, d79);
	nand (d92, d74, d77);
	xnor (d93, d68, d69);
	xnor (d94, d68, d79);
	nand (d95, d81);
	nand (d96, d79, d80);
	and (d97, d65);
	nor (d98, d65, d80);
	xor (d99, d80, d81);
	xnor (d100, d65, d73);
	or (d101, d76, d79);
	nand (d102, d72, d76);
	nand (d103, d68, d83);
	nor (d104, d69, d80);
	and (d105, d67, d83);
	nand (d106, d68, d73);
	nor (d107, d72, d81);
	nand (d108, d65, d73);
	xnor (d109, d66, d80);
	nor (d110, d66, d72);
	or (d111, d65, d71);
	buf (d112, d8);
	buf (d113, d76);
	xnor (d114, d67, d78);
	not (d115, d34);
	xnor (d116, d74, d78);
	buf (d117, d9);
	xnor (d118, d78, d79);
	and (d119, d67, d69);
	nor (d120, d70, d74);
	not (d121, d42);
	or (d122, d76, d78);
	nor (d123, d69, d78);
	xor (d124, d77);
	and (d125, d66, d68);
	buf (d126, d10);
	and (d127, d66, d74);
	not (d128, d41);
	nand (d129, d69, d76);
	nand (d130, d74, d75);
	not (d131, d75);
	xor (d132, d77, d80);
	nor (d133, d67, d78);
	nand (d134, d80, d83);
	or (d135, d67, d80);
	not (d136, d5);
	buf (d137, d44);
	nand (d138, d77, d82);
	not (d139, d59);
	nand (d140, d75, d83);
	buf (d141, d35);
	nand (d142, d67, d80);
	nor (d143, d69, d71);
	buf (d144, d48);
	or (d145, d80, d83);
	not (d146, d79);
	or (d147, d66);
	xnor (d148, d90, d140);
	not (d149, d36);
	xnor (d150, d129, d142);
	not (d151, d17);
	xnor (d152, d101, d118);
	xor (d153, d138, d139);
	nand (d154, d88, d108);
	and (d155, d117, d137);
	xnor (d156, d133, d134);
	or (d157, d140, d141);
	not (d158, d130);
	xnor (d159, d89, d126);
	xnor (d160, d111, d144);
	xnor (d161, d127, d147);
	nor (d162, d103, d119);
	or (d163, d89, d132);
	or (d164, d88, d118);
	buf (d165, d80);
	xor (d166, d89, d112);
	xnor (d167, d103, d129);
	not (d168, d94);
	xnor (d169, d125, d130);
	or (d170, d110, d139);
	xnor (d171, d87, d110);
	nand (d172, d98, d131);
	xnor (d173, d95, d120);
	and (d174, d106, d127);
	xnor (d175, d101, d114);
	or (d176, d107, d139);
	and (d177, d98, d117);
	xnor (d178, d86, d111);
	buf (d179, d138);
	xnor (d180, d92, d103);
	xnor (d181, d101, d103);
	nor (d182, d90, d142);
	or (d183, d92, d114);
	and (d184, d101, d133);
	xor (d185, d101, d122);
	not (d186, d70);
	buf (d187, d141);
	and (d188, d98, d133);
	nand (d189, d117, d135);
	and (d190, d87, d99);
	buf (d191, d17);
	nor (d192, d109, d122);
	buf (d193, d14);
	xor (d194, d89, d100);
	and (d195, d105, d109);
	xnor (d196, d110, d118);
	nor (d197, d108, d140);
	xnor (d198, d100, d142);
	or (d199, d107, d127);
	or (d200, d117, d132);
	buf (d201, d94);
	or (d202, d93, d139);
	xor (d203, d139, d143);
	nand (d204, d95, d136);
	xnor (d205, d108, d114);
	not (d206, d97);
	and (d207, d91, d95);
	not (d208, d58);
	xor (d209, d94, d123);
	and (d210, d89, d120);
	buf (d211, d82);
	buf (d212, d79);
	not (d213, d66);
	nor (d214, d96, d137);
	xnor (d215, d100, d118);
	xor (d216, d88, d130);
	and (d217, d90, d146);
	xor (d218, d160, d164);
	nand (d219, d148, d208);
	xnor (d220, d178, d200);
	or (d221, d175, d197);
	and (d222, d168, d177);
	nand (d223, d172, d190);
	not (d224, d7);
	or (d225, d158, d203);
	xnor (d226, d149, d150);
	not (d227, d43);
	nor (d228, d195, d197);
	not (d229, d13);
	not (d230, d56);
	xor (d231, d171, d207);
	nor (d232, d190, d214);
	nor (d233, d155, d210);
	not (d234, d38);
	xor (d235, d148, d186);
	or (d236, d186, d215);
	nand (d237, d169, d189);
	not (d238, d117);
	and (d239, d184, d215);
	buf (d240, d142);
	and (d241, d160, d198);
	or (d242, d164, d196);
	nand (d243, d158, d174);
	nand (d244, d149, d205);
	nand (d245, d164, d208);
	buf (d246, d115);
	buf (d247, d147);
	nor (d248, d152, d163);
	and (d249, d179, d210);
	xnor (d250, d156, d171);
	nor (d251, d185, d202);
	xor (d252, d181, d213);
	xor (d253, d187, d200);
	or (d254, d180, d185);
	buf (d255, d37);
	xor (d256, d158, d213);
	and (d257, d201, d212);
	buf (d258, d95);
	and (d259, d156, d158);
	nor (d260, d175, d213);
	not (d261, d194);
	nor (d262, d180, d205);
	nor (d263, d163, d176);
	nand (d264, d197, d213);
	or (d265, d166, d210);
	nor (d266, d224, d226);
	xor (d267, d249, d250);
	and (d268, d236, d256);
	nand (d269, d219, d228);
	not (d270, d231);
	and (d271, d260, d261);
	nand (d272, d237, d259);
	xor (d273, d231, d257);
	xor (d274, d257, d258);
	xnor (d275, d225, d244);
	buf (d276, d40);
	and (d277, d225, d258);
	not (d278, d235);
	not (d279, d170);
	or (d280, d233, d254);
	nor (d281, d240, d263);
	buf (d282, d193);
	nand (d283, d237, d238);
	not (d284, d119);
	and (d285, d255, d258);
	xor (d286, d224, d259);
	xor (d287, d252, d260);
	xor (d288, d227, d247);
	buf (d289, d258);
	nand (d290, d243, d258);
	or (d291, d235, d265);
	xor (d292, d220, d255);
	xnor (d293, d226, d254);
	nand (d294, d237, d239);
	not (d295, d160);
	xnor (d296, d224, d265);
	xor (d297, d233, d236);
	xnor (d298, d243, d256);
	not (d299, d154);
	nor (d300, d234, d263);
	xor (d301, d231, d252);
	xor (d302, d218, d228);
	xnor (d303, d249, d262);
	xnor (d304, d229, d255);
	buf (d305, d97);
	nor (d306, d235, d261);
	buf (d307, d77);
	nor (d308, d228, d258);
	xnor (d309, d231, d256);
	and (d310, d226, d262);
	nand (d311, d232, d256);
	nor (d312, d248, d265);
	not (d313, d39);
	buf (d314, d107);
	and (d315, d231, d244);
	nor (d316, d223, d230);
	buf (d317, d100);
	xnor (d318, d226, d264);
	and (d319, d229, d233);
	nor (d320, d241, d247);
	xor (d321, d220, d243);
	buf (d322, d217);
	buf (d323, d189);
	not (d324, d53);
	xor (d325, d230, d232);
	and (d326, d219, d241);
	buf (d327, d16);
	not (d328, d108);
	xor (d329, d247, d253);
	or (d330, d250, d259);
	xor (d331, d222, d234);
	xnor (d332, d241, d253);
	buf (d333, d54);
	buf (d334, d36);
	buf (d335, d111);
	nand (d336, d234, d239);
	and (d337, d220, d251);
	xnor (d338, d235, d243);
	nand (d339, d231, d235);
	buf (d340, d197);
	or (d341, d219, d261);
	not (d342, d28);
	not (d343, d152);
	nor (d344, d228, d257);
	buf (d345, d229);
	nand (d346, d226, d243);
	not (d347, d188);
	nand (d348, d219, d236);
	nand (d349, d244, d245);
	not (d350, d147);
	buf (d351, d190);
	nand (d352, d261, d264);
	xnor (d353, d244, d260);
	nor (d354, d248, d258);
	not (d355, d174);
	assign f1 = d330;
	assign f2 = d290;
	assign f3 = d313;
	assign f4 = d305;
	assign f5 = d341;
	assign f6 = d312;
	assign f7 = d316;
	assign f8 = d299;
endmodule
