module CCGRCG30( x0, x1, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17 );

	input x0, x1;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314, d315, d316, d317, d318, d319, d320, d321, d322, d323, d324, d325, d326, d327, d328, d329, d330, d331, d332, d333, d334, d335, d336, d337, d338, d339, d340, d341, d342, d343, d344, d345, d346, d347, d348, d349, d350, d351, d352, d353, d354, d355, d356, d357, d358, d359, d360, d361, d362, d363, d364, d365, d366, d367, d368, d369, d370, d371, d372, d373, d374, d375, d376, d377, d378, d379, d380, d381, d382, d383, d384, d385, d386, d387, d388, d389, d390, d391, d392, d393, d394, d395, d396, d397;

	buf (d1, x1);
	xor (d2, x1);
	buf (d3, x0);
	nor (d4, x0);
	nand (d5, x0, x1);
	and (d6, x0, x1);
	or (d7, x1);
	or (d8, x0);
	nand (d9, x0, x1);
	not (d10, x0);
	and (d11, x1);
	xor (d12, x0, x1);
	xor (d13, x0, x1);
	nand (d14, x1);
	xnor (d15, x0, x1);
	not (d16, x1);
	nor (d17, x1);
	xnor (d18, x0);
	xor (d19, x0);
	or (d20, d5, d14);
	and (d21, d7, d9);
	buf (d22, d11);
	not (d23, d3);
	xor (d24, d11, d12);
	nor (d25, d1, d4);
	nor (d26, d1, d16);
	nor (d27, d21, d25);
	and (d28, d20, d21);
	buf (d29, d3);
	xnor (d30, d23);
	and (d31, d21, d22);
	nor (d32, d21, d22);
	nor (d33, d24, d25);
	xnor (d34, d21, d25);
	not (d35, d1);
	buf (d36, d4);
	or (d37, d21, d25);
	buf (d38, d6);
	buf (d39, d18);
	nor (d40, d20, d25);
	buf (d41, d9);
	or (d42, d22, d25);
	nand (d43, d20, d23);
	xor (d44, d20, d25);
	xnor (d45, d22, d26);
	not (d46, d24);
	not (d47, d6);
	and (d48, d20, d22);
	nand (d49, d24, d26);
	nand (d50, d20, d22);
	nand (d51, d23, d24);
	buf (d52, d15);
	and (d53, d20);
	and (d54, d25);
	xnor (d55, d20, d23);
	nor (d56, d23, d24);
	not (d57, d19);
	not (d58, d21);
	not (d59, d12);
	or (d60, d21, d26);
	xor (d61, d23, d25);
	or (d62, d23, d25);
	nand (d63, d20, d22);
	or (d64, d21, d22);
	xnor (d65, d21, d23);
	xor (d66, d25);
	or (d67, d22, d26);
	and (d68, d20, d23);
	not (d69, d16);
	xnor (d70, d21, d26);
	nor (d71, d20);
	xor (d72, d21, d24);
	xnor (d73, d26);
	nand (d74, d21, d23);
	nand (d75, d20, d21);
	xor (d76, d23);
	and (d77, d25, d26);
	and (d78, d23, d24);
	nor (d79, d22, d24);
	nor (d80, d22, d25);
	and (d81, d20, d25);
	xnor (d82, d21, d24);
	nand (d83, d21, d26);
	xor (d84, d20, d25);
	not (d85, d23);
	buf (d86, d8);
	nand (d87, d21, d25);
	or (d88, d22);
	nor (d89, d24, d26);
	and (d90, d42, d76);
	buf (d91, d71);
	not (d92, d11);
	nand (d93, d60, d76);
	and (d94, d32, d52);
	not (d95, d44);
	xor (d96, d59, d64);
	xor (d97, d46, d84);
	xor (d98, d53, d60);
	buf (d99, d55);
	xnor (d100, d40, d49);
	nor (d101, d56, d68);
	nor (d102, d44, d72);
	nand (d103, d50, d84);
	or (d104, d39, d47);
	not (d105, d38);
	buf (d106, d66);
	xnor (d107, d47, d54);
	and (d108, d54);
	nor (d109, d39, d68);
	and (d110, d68, d86);
	and (d111, d37, d43);
	xnor (d112, d54, d83);
	not (d113, d9);
	nor (d114, d50, d66);
	or (d115, d68, d70);
	nor (d116, d35, d38);
	and (d117, d51, d74);
	or (d118, d42, d52);
	xnor (d119, d40, d82);
	nor (d120, d88, d89);
	and (d121, d62, d88);
	not (d122, d84);
	nand (d123, d86, d88);
	nor (d124, d68, d86);
	nand (d125, d52, d85);
	not (d126, d66);
	nor (d127, d40, d89);
	buf (d128, d40);
	buf (d129, d25);
	not (d130, d59);
	or (d131, d33, d43);
	nand (d132, d45, d84);
	xnor (d133, d60, d66);
	nor (d134, d67, d76);
	and (d135, d51, d61);
	not (d136, d8);
	buf (d137, d85);
	nor (d138, d46);
	nor (d139, d86, d88);
	nand (d140, d47, d75);
	or (d141, d36, d83);
	nand (d142, d31, d89);
	xnor (d143, d34, d80);
	or (d144, d35, d49);
	or (d145, d72);
	nor (d146, d29, d75);
	and (d147, d59, d75);
	or (d148, d104, d112);
	nand (d149, d93, d123);
	buf (d150, d56);
	or (d151, d100, d145);
	xor (d152, d120);
	or (d153, d92, d117);
	and (d154, d90, d134);
	not (d155, d49);
	nor (d156, d102, d103);
	nor (d157, d120, d125);
	nand (d158, d95, d102);
	xor (d159, d116, d141);
	xnor (d160, d100, d132);
	buf (d161, d93);
	nand (d162, d95, d107);
	and (d163, d128, d134);
	nor (d164, d92, d114);
	buf (d165, d147);
	nand (d166, d92, d113);
	xnor (d167, d105, d112);
	and (d168, d108, d132);
	or (d169, d93, d119);
	nor (d170, d109, d117);
	or (d171, d119, d139);
	buf (d172, d60);
	and (d173, d103, d147);
	xnor (d174, d121, d146);
	buf (d175, d80);
	buf (d176, d50);
	xnor (d177, d109, d138);
	nand (d178, d105, d110);
	xor (d179, d93, d114);
	or (d180, d95, d132);
	xor (d181, d146, d147);
	and (d182, d99, d141);
	or (d183, d98, d122);
	xor (d184, d101, d138);
	nand (d185, d111, d136);
	and (d186, d90, d136);
	not (d187, d41);
	nor (d188, d91, d93);
	or (d189, d92, d115);
	nor (d190, d100, d110);
	and (d191, d105, d136);
	or (d192, d152, d165);
	xor (d193, d163, d168);
	and (d194, d152, d184);
	and (d195, d155, d188);
	nor (d196, d167, d177);
	or (d197, d148, d190);
	nand (d198, d165, d170);
	and (d199, d154, d162);
	xnor (d200, d150, d189);
	xor (d201, d152, d186);
	xnor (d202, d172, d180);
	nand (d203, d161, d178);
	or (d204, d157, d170);
	or (d205, d156, d157);
	xor (d206, d153, d172);
	xnor (d207, d167, d179);
	not (d208, d69);
	xnor (d209, d183, d185);
	nor (d210, d151, d165);
	nand (d211, d164);
	not (d212, d177);
	xnor (d213, d159, d162);
	buf (d214, d110);
	or (d215, d152, d181);
	xor (d216, d155, d162);
	buf (d217, d122);
	nor (d218, d163, d168);
	buf (d219, d30);
	xnor (d220, d163, d189);
	and (d221, d162, d175);
	buf (d222, d74);
	not (d223, d143);
	xor (d224, d169, d190);
	not (d225, d62);
	nand (d226, d178, d188);
	and (d227, d177, d186);
	buf (d228, d20);
	nand (d229, d151, d164);
	and (d230, d162, d185);
	nor (d231, d150, d151);
	nand (d232, d171, d177);
	xor (d233, d148, d168);
	nand (d234, d148, d186);
	or (d235, d162, d178);
	not (d236, d51);
	nand (d237, d176, d180);
	not (d238, d99);
	or (d239, d154, d180);
	buf (d240, d96);
	or (d241, d157, d177);
	xor (d242, d158, d160);
	nor (d243, d163, d183);
	not (d244, d128);
	or (d245, d184);
	or (d246, d153, d160);
	nor (d247, d170, d187);
	or (d248, d152, d159);
	not (d249, d83);
	buf (d250, d126);
	nand (d251, d182, d188);
	or (d252, d168, d186);
	nor (d253, d159, d190);
	not (d254, d150);
	xnor (d255, d160, d171);
	xnor (d256, d154, d182);
	buf (d257, d91);
	xnor (d258, d205, d242);
	nor (d259, d218, d255);
	nand (d260, d211, d223);
	not (d261, d159);
	not (d262, d232);
	xor (d263, d192, d240);
	or (d264, d193, d231);
	nor (d265, d195, d227);
	xor (d266, d215, d226);
	not (d267, d81);
	xnor (d268, d218, d238);
	and (d269, d195, d250);
	or (d270, d221, d246);
	nor (d271, d207, d217);
	nand (d272, d216, d237);
	buf (d273, d94);
	nand (d274, d222, d236);
	buf (d275, d136);
	and (d276, d213, d231);
	nor (d277, d207, d255);
	and (d278, d225, d226);
	and (d279, d198);
	not (d280, d78);
	xnor (d281, d222, d252);
	xnor (d282, d195, d214);
	xor (d283, d226, d250);
	nand (d284, d192, d195);
	not (d285, d97);
	nor (d286, d203, d226);
	nor (d287, d207, d243);
	nor (d288, d207, d247);
	buf (d289, d123);
	xnor (d290, d202, d244);
	not (d291, d18);
	not (d292, d241);
	nand (d293, d196, d230);
	xnor (d294, d228, d244);
	not (d295, d39);
	xnor (d296, d243, d247);
	or (d297, d199, d201);
	or (d298, d200, d245);
	nand (d299, d197, d240);
	not (d300, d122);
	buf (d301, d98);
	not (d302, d17);
	and (d303, d219, d228);
	nor (d304, d217, d238);
	nand (d305, d199, d206);
	xnor (d306, d207, d209);
	buf (d307, d35);
	or (d308, d196, d243);
	not (d309, d104);
	xor (d310, d199, d243);
	nor (d311, d192, d248);
	xnor (d312, d233, d245);
	not (d313, d186);
	nor (d314, d216, d233);
	xnor (d315, d203, d227);
	not (d316, d219);
	nand (d317, d217, d254);
	or (d318, d201, d249);
	nand (d319, d222, d237);
	not (d320, d142);
	not (d321, d71);
	xor (d322, d204, d209);
	and (d323, d228, d229);
	and (d324, d234, d252);
	xor (d325, d247, d250);
	nor (d326, d201, d226);
	or (d327, d220, d244);
	xor (d328, d198, d246);
	nor (d329, d192, d217);
	xnor (d330, d195, d200);
	buf (d331, d51);
	nor (d332, d208, d244);
	nand (d333, d240, d250);
	or (d334, d193, d208);
	buf (d335, d101);
	and (d336, d217, d231);
	xor (d337, d213, d245);
	xnor (d338, d203, d247);
	nand (d339, d206, d234);
	nand (d340, d213, d219);
	not (d341, d222);
	xor (d342, d220, d246);
	nor (d343, d201, d222);
	buf (d344, d124);
	nand (d345, d330, d335);
	xnor (d346, d259, d290);
	xor (d347, d312, d323);
	nor (d348, d292, d318);
	nand (d349, d266, d293);
	nand (d350, d263, d339);
	and (d351, d270, d292);
	or (d352, d281, d307);
	or (d353, d296, d330);
	or (d354, d302, d344);
	and (d355, d330, d339);
	nor (d356, d258, d280);
	not (d357, d147);
	xnor (d358, d259, d314);
	nand (d359, d293, d329);
	xor (d360, d279, d337);
	or (d361, d260, d317);
	nand (d362, d283, d322);
	not (d363, d290);
	nand (d364, d260, d341);
	nand (d365, d297, d330);
	not (d366, d326);
	xnor (d367, d282, d337);
	nand (d368, d284, d297);
	buf (d369, d262);
	nor (d370, d271, d292);
	xnor (d371, d276, d304);
	buf (d372, d250);
	or (d373, d280, d306);
	xnor (d374, d273, d342);
	nand (d375, d308, d334);
	nor (d376, d263, d308);
	nand (d377, d305, d314);
	xor (d378, d258, d319);
	nand (d379, d270, d278);
	or (d380, d290, d292);
	nor (d381, d277, d311);
	not (d382, d255);
	buf (d383, d302);
	buf (d384, d81);
	or (d385, d266, d308);
	nor (d386, d291);
	nand (d387, d257, d304);
	not (d388, d70);
	and (d389, d321, d341);
	or (d390, d338, d344);
	nand (d391, d314, d337);
	nand (d392, d289, d333);
	and (d393, d309, d343);
	nand (d394, d325, d341);
	not (d395, d315);
	not (d396, d251);
	xnor (d397, d267, d319);
	assign f1 = d382;
	assign f2 = d361;
	assign f3 = d387;
	assign f4 = d345;
	assign f5 = d377;
	assign f6 = d379;
	assign f7 = d379;
	assign f8 = d396;
	assign f9 = d387;
	assign f10 = d367;
	assign f11 = d387;
	assign f12 = d391;
	assign f13 = d368;
	assign f14 = d378;
	assign f15 = d355;
	assign f16 = d357;
	assign f17 = d387;
endmodule
