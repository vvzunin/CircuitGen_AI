module CCGRCG43( x0, x1, x2, f1, f2, f3, f4 );

	input x0, x1, x2;
	output f1, f2, f3, f4;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314, d315, d316, d317, d318, d319, d320, d321, d322, d323, d324, d325, d326, d327, d328, d329, d330, d331, d332, d333, d334, d335, d336, d337, d338, d339, d340, d341, d342, d343, d344, d345, d346, d347, d348, d349, d350, d351, d352, d353, d354, d355, d356, d357, d358, d359, d360, d361, d362, d363, d364, d365, d366, d367, d368, d369, d370, d371, d372, d373, d374, d375, d376, d377, d378, d379, d380, d381, d382, d383, d384, d385, d386, d387, d388, d389, d390, d391, d392, d393, d394, d395, d396, d397, d398, d399, d400, d401, d402, d403, d404, d405, d406, d407, d408, d409, d410, d411, d412, d413, d414, d415, d416, d417, d418, d419, d420, d421, d422, d423, d424, d425, d426, d427, d428, d429, d430, d431, d432, d433, d434, d435, d436, d437, d438, d439, d440, d441, d442, d443, d444, d445, d446, d447, d448, d449, d450, d451, d452, d453, d454, d455, d456, d457, d458, d459, d460, d461, d462, d463, d464, d465, d466, d467, d468, d469, d470, d471, d472, d473, d474, d475, d476, d477, d478, d479, d480, d481, d482, d483, d484, d485, d486, d487, d488, d489, d490, d491, d492, d493, d494, d495, d496, d497, d498, d499, d500, d501, d502, d503, d504, d505, d506, d507, d508, d509, d510, d511, d512, d513, d514, d515, d516, d517, d518, d519, d520, d521, d522, d523, d524, d525, d526, d527, d528, d529, d530, d531, d532, d533, d534, d535, d536, d537, d538, d539, d540, d541, d542, d543, d544, d545, d546, d547, d548, d549, d550, d551, d552, d553, d554, d555, d556;

	nand (d1, x0, x2);
	and (d2, x2);
	xor (d3, x1, x2);
	xnor (d4, x1, x2);
	or (d5, x1);
	not (d6, x2);
	buf (d7, x2);
	xnor (d8, x0);
	xor (d9, x1);
	or (d10, x0, x2);
	or (d11, x1, x2);
	nor (d12, x1, x2);
	xor (d13, x0, x1);
	not (d14, x0);
	xnor (d15, x1);
	xor (d16, x0, x2);
	nand (d17, x1, x2);
	nand (d18, x0);
	xor (d19, x0);
	xnor (d20, x0, x2);
	xor (d21, x0, x2);
	nand (d22, x1);
	or (d23, x0, x1);
	buf (d24, x0);
	xor (d25, x1, x2);
	or (d26, x2);
	nand (d27, x0, x1);
	and (d28, x0, x2);
	and (d29, x1);
	buf (d30, x1);
	not (d31, x1);
	nor (d32, x0, x1);
	nand (d33, x2);
	or (d34, x1, x2);
	nand (d35, x1, x2);
	xor (d36, x2);
	xor (d37, x0, x1);
	nor (d38, x1, x2);
	and (d39, x1, x2);
	or (d40, x0);
	or (d41, x0, x2);
	nor (d42, x0, x2);
	nor (d43, x1);
	and (d44, x0);
	or (d45, x0, x1);
	and (d46, x0, x2);
	xnor (d47, x2);
	and (d48, x0, x1);
	xnor (d49, x0, x1);
	xnor (d50, d16, d24);
	and (d51, d2, d19);
	xor (d52, d29, d42);
	and (d53, d11, d18);
	buf (d54, d28);
	not (d55, d39);
	not (d56, d22);
	nor (d57, d5, d48);
	nor (d58, d7, d20);
	or (d59, d4, d47);
	or (d60, d3, d38);
	and (d61, d5, d48);
	or (d62, d5, d27);
	or (d63, d4, d20);
	not (d64, d35);
	xor (d65, d39, d45);
	nand (d66, d21, d43);
	and (d67, d7, d11);
	or (d68, d17, d46);
	not (d69, d46);
	xor (d70, d55, d57);
	nor (d71, d62, d63);
	or (d72, d52, d61);
	xnor (d73, d57, d61);
	and (d74, d54, d59);
	and (d75, d53, d63);
	xnor (d76, d50);
	nand (d77, d51, d61);
	nand (d78, d51, d60);
	not (d79, d24);
	and (d80, d52, d62);
	not (d81, d44);
	and (d82, d54, d56);
	nand (d83, d53, d54);
	nand (d84, d53, d56);
	nor (d85, d60, d65);
	nand (d86, d61, d62);
	not (d87, d28);
	nand (d88, d51, d53);
	xor (d89, d60, d65);
	nor (d90, d59, d65);
	xor (d91, d50, d60);
	xnor (d92, d57, d67);
	not (d93, d30);
	buf (d94, d40);
	not (d95, d27);
	not (d96, d19);
	nand (d97, d52, d61);
	nor (d98, d55, d56);
	nor (d99, d51, d60);
	xor (d100, d54, d65);
	nor (d101, d66, d68);
	and (d102, d54, d58);
	or (d103, d60, d65);
	xnor (d104, d56, d61);
	nand (d105, d57, d67);
	xnor (d106, d52, d65);
	or (d107, d56, d63);
	xor (d108, d50, d64);
	xor (d109, d51, d54);
	or (d110, d57, d58);
	or (d111, d63, d68);
	nand (d112, d51, d64);
	buf (d113, d8);
	and (d114, d52, d65);
	xnor (d115, d51, d62);
	or (d116, d52, d53);
	not (d117, d47);
	and (d118, d57, d65);
	buf (d119, d66);
	nor (d120, d57, d68);
	nor (d121, d53, d63);
	not (d122, d12);
	xnor (d123, d63);
	xnor (d124, d52, d68);
	not (d125, d67);
	nand (d126, d57, d65);
	xor (d127, d61);
	and (d128, d56, d67);
	or (d129, d64, d66);
	or (d130, d56, d65);
	nor (d131, d55, d68);
	nand (d132, d51, d67);
	nor (d133, d52, d53);
	buf (d134, d63);
	xor (d135, d50, d62);
	and (d136, d53, d59);
	or (d137, d68);
	xor (d138, d57, d67);
	or (d139, d58, d66);
	xnor (d140, d50, d57);
	and (d141, d58, d59);
	or (d142, d53, d55);
	xor (d143, d55, d68);
	and (d144, d56, d60);
	and (d145, d90);
	or (d146, d113, d116);
	buf (d147, d23);
	or (d148, d99, d116);
	xor (d149, d74, d137);
	nand (d150, d112, d137);
	and (d151, d77, d98);
	nand (d152, d88, d95);
	not (d153, d8);
	nor (d154, d76, d105);
	and (d155, d113, d132);
	nor (d156, d86, d122);
	nor (d157, d78, d108);
	xor (d158, d100, d120);
	nor (d159, d92, d132);
	buf (d160, d140);
	not (d161, d83);
	nor (d162, d80, d125);
	xor (d163, d71, d101);
	xnor (d164, d90, d111);
	nand (d165, d86, d114);
	nand (d166, d73, d92);
	xnor (d167, d69, d110);
	nand (d168, d75, d133);
	xor (d169, d69, d72);
	xnor (d170, d131, d134);
	nor (d171, d70, d92);
	buf (d172, d143);
	nand (d173, d69, d87);
	nand (d174, d82, d122);
	xnor (d175, d70);
	or (d176, d99, d120);
	not (d177, d124);
	nor (d178, d95, d108);
	nand (d179, d98, d139);
	xnor (d180, d87, d89);
	and (d181, d159, d172);
	xor (d182, d167);
	buf (d183, d18);
	nand (d184, d147, d169);
	nand (d185, d145, d147);
	xor (d186, d160, d161);
	or (d187, d164, d176);
	xnor (d188, d151, d167);
	not (d189, d76);
	buf (d190, d74);
	xnor (d191, d157, d158);
	xnor (d192, d152, d174);
	not (d193, d162);
	or (d194, d164, d178);
	xor (d195, d145, d152);
	buf (d196, d110);
	and (d197, d146, d180);
	xnor (d198, d147, d179);
	nand (d199, d163, d171);
	nand (d200, d149, d162);
	buf (d201, d121);
	xnor (d202, d153, d157);
	buf (d203, d115);
	or (d204, d147, d161);
	nor (d205, d152, d170);
	or (d206, d165, d170);
	xnor (d207, d147, d177);
	xor (d208, d154, d172);
	xnor (d209, d167, d177);
	or (d210, d175, d176);
	xnor (d211, d147, d167);
	or (d212, d146, d159);
	xor (d213, d168, d169);
	nand (d214, d150, d160);
	and (d215, d171);
	nor (d216, d145, d163);
	or (d217, d150, d153);
	xnor (d218, d161, d171);
	and (d219, d161, d179);
	nor (d220, d162, d169);
	nor (d221, d167, d173);
	nor (d222, d164, d173);
	or (d223, d152, d159);
	or (d224, d151, d167);
	nand (d225, d147, d170);
	and (d226, d167);
	nand (d227, d160, d169);
	xnor (d228, d156, d163);
	nor (d229, d146, d153);
	or (d230, d164, d169);
	xnor (d231, d155, d179);
	xor (d232, d161, d166);
	or (d233, d165, d170);
	and (d234, d175, d177);
	nand (d235, d148, d178);
	buf (d236, d173);
	xnor (d237, d159, d175);
	buf (d238, d137);
	and (d239, d170, d171);
	xnor (d240, d151, d172);
	nand (d241, d156, d171);
	nand (d242, d175);
	xnor (d243, d153, d178);
	or (d244, d164, d167);
	nand (d245, d179, d180);
	xor (d246, d166, d178);
	or (d247, d146, d178);
	nor (d248, d156, d177);
	xnor (d249, d151, d153);
	nor (d250, d147, d164);
	buf (d251, d96);
	and (d252, d168, d179);
	or (d253, d154, d177);
	and (d254, d168, d175);
	or (d255, d148, d166);
	or (d256, d151, d153);
	nand (d257, d157, d179);
	and (d258, d160, d165);
	nor (d259, d177, d179);
	xnor (d260, d145, d146);
	xor (d261, d147, d160);
	and (d262, d151, d167);
	buf (d263, d154);
	nor (d264, d149, d157);
	xor (d265, d152, d174);
	xor (d266, d152, d160);
	nor (d267, d157, d174);
	xor (d268, d157, d173);
	not (d269, d53);
	or (d270, d150, d159);
	nor (d271, d151, d173);
	nor (d272, d145, d169);
	or (d273, d159, d171);
	nor (d274, d155, d164);
	not (d275, d267);
	xnor (d276, d221, d224);
	nand (d277, d206, d260);
	and (d278, d214, d255);
	nor (d279, d201, d265);
	not (d280, d180);
	and (d281, d197, d270);
	nor (d282, d212, d250);
	buf (d283, d93);
	nor (d284, d194, d215);
	nand (d285, d224, d252);
	or (d286, d217, d249);
	xnor (d287, d202, d233);
	xor (d288, d232, d249);
	not (d289, d32);
	and (d290, d231, d248);
	nor (d291, d183, d197);
	nor (d292, d210, d216);
	xnor (d293, d191, d274);
	xor (d294, d236, d270);
	not (d295, d62);
	nor (d296, d183, d219);
	nand (d297, d209, d265);
	buf (d298, d142);
	xnor (d299, d204, d207);
	not (d300, d183);
	nand (d301, d251, d265);
	or (d302, d246, d250);
	or (d303, d252, d253);
	xor (d304, d205, d229);
	buf (d305, d57);
	not (d306, d222);
	and (d307, d181, d254);
	nand (d308, d195, d212);
	buf (d309, d111);
	xnor (d310, d252, d274);
	nor (d311, d254, d274);
	buf (d312, d10);
	xnor (d313, d211, d266);
	xor (d314, d195, d201);
	and (d315, d249, d259);
	xor (d316, d234, d252);
	buf (d317, d109);
	or (d318, d220, d238);
	xnor (d319, d208, d241);
	and (d320, d181, d221);
	or (d321, d218, d260);
	and (d322, d191, d210);
	xnor (d323, d191, d215);
	or (d324, d190, d228);
	or (d325, d198, d237);
	or (d326, d183, d261);
	xnor (d327, d186, d211);
	and (d328, d204, d246);
	xor (d329, d220, d268);
	nand (d330, d244, d253);
	or (d331, d186, d246);
	buf (d332, d266);
	nor (d333, d222, d244);
	not (d334, d188);
	nand (d335, d185, d250);
	not (d336, d172);
	and (d337, d187, d240);
	and (d338, d286, d315);
	and (d339, d280, d325);
	nor (d340, d292, d308);
	and (d341, d317, d318);
	and (d342, d295, d300);
	nor (d343, d292, d321);
	and (d344, d293, d296);
	not (d345, d168);
	not (d346, d310);
	and (d347, d280, d307);
	or (d348, d301, d321);
	buf (d349, d208);
	nor (d350, d309, d335);
	xnor (d351, d293, d300);
	xor (d352, d281, d329);
	nand (d353, d295, d299);
	not (d354, d224);
	and (d355, d307, d322);
	or (d356, d305, d332);
	xor (d357, d289, d295);
	xnor (d358, d277, d286);
	nor (d359, d289, d315);
	or (d360, d297, d337);
	not (d361, d181);
	xnor (d362, d280, d323);
	buf (d363, d67);
	xnor (d364, d317, d324);
	or (d365, d298, d323);
	and (d366, d298, d308);
	xnor (d367, d281, d326);
	and (d368, d303, d328);
	nor (d369, d293, d306);
	xnor (d370, d284, d297);
	nor (d371, d296, d333);
	or (d372, d281, d304);
	xor (d373, d280, d297);
	nand (d374, d279, d328);
	not (d375, d217);
	xnor (d376, d325, d337);
	xor (d377, d288, d309);
	nor (d378, d315, d318);
	xor (d379, d325, d331);
	or (d380, d300, d311);
	and (d381, d278, d325);
	and (d382, d281, d283);
	xor (d383, d289, d310);
	nand (d384, d278, d299);
	buf (d385, d302);
	or (d386, d276, d316);
	xnor (d387, d278, d289);
	buf (d388, d100);
	xnor (d389, d296, d303);
	and (d390, d299, d326);
	or (d391, d281, d290);
	nand (d392, d300, d308);
	nand (d393, d285, d331);
	and (d394, d280, d332);
	buf (d395, d310);
	and (d396, d338, d372);
	xnor (d397, d370, d385);
	or (d398, d357, d360);
	nand (d399, d358, d365);
	nand (d400, d351, d354);
	and (d401, d341, d342);
	nor (d402, d350, d382);
	and (d403, d341, d383);
	not (d404, d137);
	buf (d405, d257);
	nor (d406, d379, d391);
	buf (d407, d159);
	xnor (d408, d340, d344);
	nor (d409, d379, d386);
	or (d410, d355, d375);
	xnor (d411, d369, d392);
	nand (d412, d362, d369);
	xor (d413, d362, d373);
	or (d414, d359, d363);
	nand (d415, d356, d388);
	nand (d416, d340, d360);
	or (d417, d347, d350);
	nand (d418, d341, d391);
	buf (d419, d294);
	buf (d420, d144);
	buf (d421, d24);
	buf (d422, d242);
	nor (d423, d352, d392);
	or (d424, d350, d359);
	and (d425, d340, d346);
	xor (d426, d390, d395);
	not (d427, d231);
	xor (d428, d345, d387);
	nand (d429, d356, d361);
	nand (d430, d384, d388);
	and (d431, d340, d379);
	nor (d432, d356, d376);
	nor (d433, d355, d364);
	nor (d434, d369, d377);
	nand (d435, d382, d392);
	xor (d436, d342, d387);
	nor (d437, d353, d375);
	buf (d438, d315);
	or (d439, d342, d348);
	xor (d440, d342, d392);
	nand (d441, d364, d386);
	xor (d442, d341, d387);
	nor (d443, d378, d387);
	not (d444, d147);
	nor (d445, d345, d359);
	buf (d446, d47);
	nand (d447, d370, d386);
	not (d448, d171);
	or (d449, d389, d391);
	not (d450, d292);
	xor (d451, d354, d374);
	or (d452, d351, d391);
	not (d453, d153);
	buf (d454, d324);
	nor (d455, d357, d386);
	xnor (d456, d369, d382);
	xor (d457, d345, d384);
	and (d458, d342, d373);
	not (d459, d107);
	nand (d460, d343, d387);
	xor (d461, d373, d378);
	buf (d462, d12);
	nor (d463, d363, d385);
	xor (d464, d364, d382);
	xnor (d465, d348, d375);
	nand (d466, d356, d392);
	xor (d467, d368, d377);
	nand (d468, d361, d379);
	xnor (d469, d378, d384);
	or (d470, d377, d388);
	xnor (d471, d377, d390);
	or (d472, d380, d394);
	nor (d473, d356, d385);
	nor (d474, d348, d386);
	nor (d475, d390, d391);
	xnor (d476, d368, d376);
	nor (d477, d344, d351);
	or (d478, d350, d361);
	nor (d479, d358, d374);
	xor (d480, d350, d392);
	and (d481, d349, d371);
	buf (d482, d41);
	nor (d483, d358, d380);
	xor (d484, d367, d381);
	and (d485, d357, d378);
	nand (d486, d343, d383);
	buf (d487, d87);
	not (d488, d302);
	or (d489, d467, d473);
	not (d490, d48);
	or (d491, d461, d464);
	buf (d492, d102);
	xor (d493, d444, d474);
	xor (d494, d454, d471);
	xor (d495, d424, d437);
	not (d496, d254);
	xnor (d497, d409, d459);
	not (d498, d210);
	or (d499, d402, d423);
	xor (d500, d433, d456);
	nand (d501, d460, d479);
	xnor (d502, d452, d469);
	or (d503, d413, d445);
	nor (d504, d414, d462);
	xnor (d505, d471, d484);
	nor (d506, d406, d486);
	or (d507, d445, d475);
	nand (d508, d449, d473);
	or (d509, d402, d467);
	nand (d510, d399, d442);
	not (d511, d470);
	buf (d512, d58);
	and (d513, d432, d434);
	xnor (d514, d450, d474);
	xnor (d515, d396, d410);
	or (d516, d428, d434);
	not (d517, d475);
	not (d518, d298);
	or (d519, d430, d479);
	xnor (d520, d475, d483);
	xnor (d521, d438, d484);
	buf (d522, d367);
	and (d523, d429, d475);
	xnor (d524, d424, d450);
	not (d525, d173);
	and (d526, d399, d411);
	nor (d527, d449, d464);
	or (d528, d417, d436);
	and (d529, d453, d466);
	buf (d530, d422);
	or (d531, d446, d448);
	nand (d532, d408, d423);
	not (d533, d57);
	xnor (d534, d434, d469);
	xnor (d535, d421, d464);
	xnor (d536, d427, d472);
	not (d537, d309);
	xnor (d538, d440, d467);
	xor (d539, d453, d461);
	xor (d540, d451, d460);
	or (d541, d406, d413);
	not (d542, d319);
	not (d543, d233);
	buf (d544, d420);
	nand (d545, d451, d477);
	not (d546, d387);
	nor (d547, d437, d440);
	xnor (d548, d401, d486);
	or (d549, d441, d476);
	and (d550, d435, d448);
	or (d551, d452, d455);
	nor (d552, d470);
	and (d553, d406, d477);
	buf (d554, d423);
	and (d555, d475, d480);
	buf (d556, d198);
	assign f1 = d538;
	assign f2 = d555;
	assign f3 = d540;
	assign f4 = d518;
endmodule
