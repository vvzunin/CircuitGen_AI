module CCGRCG139( x0, x1, x2, x3, x4, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14 );

	input x0, x1, x2, x3, x4;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87;

	and (d1, x3, x4);
	or (d2, x1, x3);
	xnor (d3, x1, x4);
	xor (d4, x1, x4);
	and (d5, x1, x2);
	nor (d6, x1, x2);
	and (d7, x1, x4);
	not (d8, x1);
	nor (d9, x1, x4);
	nor (d10, x2, x4);
	or (d11, x1, x2);
	or (d12, x0, x1);
	nand (d13, x3, x4);
	nor (d14, x0, x2);
	buf (d15, x0);
	xnor (d16, x1, x2);
	nand (d17, x2);
	xnor (d18, x0);
	xor (d19, x2, x3);
	not (d20, x4);
	xnor (d21, x0, x2);
	or (d22, x0, x4);
	nand (d23, x2, x3);
	and (d24, x3);
	and (d25, x0, x1);
	and (d26, x4);
	xor (d27, x0);
	nand (d28, x0, x2);
	nand (d29, x2, x4);
	xor (d30, x0, x4);
	nor (d31, x1, x4);
	xor (d32, x3);
	or (d33, x1, x3);
	not (d34, x2);
	nor (d35, x4);
	nor (d36, x0, x3);
	nor (d37, x1, x3);
	xor (d38, x4);
	xor (d39, x1, x3);
	and (d40, x0, x3);
	or (d41, d14, d28);
	nor (d42, d9, d38);
	nor (d43, d7, d35);
	xnor (d44, d8, d30);
	nand (d45, d11, d31);
	nand (d46, d28, d31);
	or (d47, d23, d31);
	and (d48, d26, d27);
	not (d49, d26);
	xnor (d50, d15, d26);
	or (d51, d6, d33);
	and (d52, d12, d30);
	buf (d53, d11);
	or (d54, d6, d34);
	xor (d55, d23, d27);
	buf (d56, d26);
	xnor (d57, d34, d36);
	or (d58, d5, d18);
	not (d59, d33);
	xor (d60, d7, d38);
	or (d61, d15, d40);
	xnor (d62, d6, d25);
	xnor (d63, d10, d30);
	and (d64, d8, d17);
	and (d65, d17, d40);
	buf (d66, d1);
	nand (d67, d34, d35);
	xnor (d68, d5, d22);
	not (d69, d23);
	or (d70, d10, d18);
	not (d71, d25);
	or (d72, d28, d40);
	nand (d73, d18, d22);
	nand (d74, d31, d38);
	buf (d75, d36);
	and (d76, d14, d24);
	nor (d77, d7, d29);
	and (d78, d24, d32);
	nand (d79, d15, d16);
	xor (d80, d21, d22);
	xnor (d81, d10, d20);
	not (d82, d12);
	not (d83, d8);
	or (d84, d3, d32);
	xnor (d85, d26, d29);
	buf (d86, d20);
	nor (d87, d19, d36);
	assign f1 = d77;
	assign f2 = d42;
	assign f3 = d82;
	assign f4 = d62;
	assign f5 = d85;
	assign f6 = d64;
	assign f7 = d60;
	assign f8 = d77;
	assign f9 = d83;
	assign f10 = d56;
	assign f11 = d73;
	assign f12 = d45;
	assign f13 = d83;
	assign f14 = d42;
endmodule
