module CCGRCG86( x0, x1, x2, x3, f1, f2, f3, f4, f5, f6, f7 );

	input x0, x1, x2, x3;
	output f1, f2, f3, f4, f5, f6, f7;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294;

	nor (d1, x1);
	nand (d2, x1, x3);
	or (d3, x2);
	not (d4, x1);
	xor (d5, x1, x2);
	and (d6, x1, x2);
	and (d7, x1, x3);
	buf (d8, x2);
	nand (d9, x0);
	nand (d10, x1, x2);
	or (d11, x0, x3);
	not (d12, x0);
	xnor (d13, x2);
	xnor (d14, x1, x3);
	nand (d15, x2, x3);
	buf (d16, x3);
	buf (d17, x1);
	or (d18, x0, x3);
	and (d19, x2, x3);
	not (d20, x2);
	and (d21, x0, x1);
	xnor (d22, x1, x2);
	or (d23, x0, x1);
	xnor (d24, x2, x3);
	nand (d25, d3, d20);
	xnor (d26, d14, d15);
	nand (d27, d12, d19);
	xor (d28, d9, d16);
	or (d29, d9, d21);
	buf (d30, d2);
	nand (d31, d9, d15);
	not (d32, d9);
	nand (d33, d16, d19);
	and (d34, d17, d23);
	or (d35, d8, d12);
	nand (d36, d4, d8);
	nor (d37, d3, d5);
	xor (d38, d19, d21);
	not (d39, d2);
	xnor (d40, d11, d19);
	or (d41, d6, d12);
	buf (d42, d3);
	not (d43, d11);
	not (d44, d1);
	xor (d45, d9, d20);
	and (d46, d11, d15);
	or (d47, d12, d17);
	and (d48, d5, d15);
	not (d49, d16);
	or (d50, d7, d8);
	nor (d51, d4, d19);
	and (d52, d5, d18);
	not (d53, d14);
	nor (d54, d17);
	or (d55, d4, d22);
	not (d56, d15);
	and (d57, d6, d24);
	or (d58, d11, d12);
	buf (d59, d24);
	xnor (d60, d8, d10);
	nand (d61, d13, d14);
	nand (d62, d24);
	or (d63, d16, d17);
	not (d64, d6);
	nand (d65, d10, d22);
	nor (d66, d3, d9);
	nor (d67, d1, d17);
	and (d68, d13, d14);
	not (d69, d20);
	not (d70, x3);
	and (d71, d11, d14);
	nor (d72, d11, d24);
	xnor (d73, d7, d21);
	buf (d74, d13);
	xor (d75, d3, d15);
	nand (d76, d8, d11);
	or (d77, d8, d14);
	or (d78, d3, d13);
	xor (d79, d3, d9);
	xor (d80, d5, d10);
	nand (d81, d16, d21);
	nor (d82, d1, d3);
	nand (d83, d21);
	not (d84, d10);
	and (d85, d3);
	xor (d86, d13, d17);
	buf (d87, d14);
	and (d88, d2, d11);
	xnor (d89, d12, d15);
	xor (d90, d10, d18);
	or (d91, d19, d23);
	and (d92, d7, d10);
	xnor (d93, d19);
	or (d94, d4, d7);
	nor (d95, d4, d11);
	and (d96, d10, d12);
	xnor (d97, d6, d16);
	nor (d98, d4, d15);
	nor (d99, d20);
	not (d100, d13);
	nor (d101, d59, d100);
	buf (d102, d34);
	nor (d103, d64, d95);
	xor (d104, d37, d75);
	and (d105, d46, d72);
	and (d106, d32, d61);
	buf (d107, d23);
	xnor (d108, d29, d38);
	or (d109, d70, d88);
	buf (d110, d96);
	xnor (d111, d55, d86);
	nor (d112, d29, d53);
	or (d113, d48, d65);
	nor (d114, d59, d75);
	and (d115, d27, d75);
	nor (d116, d75, d90);
	xnor (d117, d74, d94);
	xor (d118, d82, d98);
	nor (d119, d39, d69);
	nor (d120, d76, d78);
	not (d121, d44);
	nand (d122, d60, d86);
	or (d123, d54, d99);
	xor (d124, d62, d95);
	not (d125, d46);
	not (d126, d8);
	nand (d127, d30, d77);
	xor (d128, d86, d88);
	buf (d129, d30);
	xor (d130, d88);
	nand (d131, d49, d62);
	and (d132, d62, d70);
	nand (d133, d34, d87);
	nand (d134, d34, d78);
	buf (d135, d16);
	buf (d136, d93);
	xnor (d137, d35, d84);
	or (d138, d28, d58);
	xnor (d139, d40, d86);
	buf (d140, d20);
	nor (d141, d32, d97);
	nor (d142, d82, d88);
	or (d143, d33, d73);
	xor (d144, d57, d99);
	and (d145, d45, d69);
	xor (d146, d76, d91);
	and (d147, d26, d83);
	not (d148, d45);
	xor (d149, d30, d43);
	xor (d150, d105, d141);
	xnor (d151, d101, d132);
	xor (d152, d105, d136);
	and (d153, d144, d149);
	xor (d154, d106, d110);
	not (d155, d42);
	or (d156, d106, d119);
	xnor (d157, d107, d146);
	xnor (d158, d136, d139);
	xor (d159, d133, d147);
	buf (d160, d105);
	and (d161, d105, d109);
	xnor (d162, d110, d143);
	nor (d163, d131, d142);
	buf (d164, d79);
	not (d165, d142);
	nor (d166, d102, d116);
	nor (d167, d101, d129);
	not (d168, d104);
	not (d169, d33);
	nand (d170, d129, d140);
	buf (d171, d67);
	buf (d172, d104);
	not (d173, d19);
	buf (d174, d48);
	nor (d175, d113, d125);
	xnor (d176, d108, d120);
	nor (d177, d123, d133);
	nor (d178, d104, d113);
	xor (d179, d129, d140);
	or (d180, d106, d149);
	nor (d181, d106, d149);
	and (d182, d119, d142);
	xnor (d183, d139);
	or (d184, d106, d145);
	buf (d185, d37);
	not (d186, d109);
	and (d187, d118, d140);
	nand (d188, d101, d106);
	buf (d189, d110);
	and (d190, d180, d188);
	nor (d191, d165, d173);
	not (d192, d151);
	nand (d193, d168, d170);
	or (d194, d160, d164);
	xor (d195, d177, d183);
	nand (d196, d154, d178);
	xnor (d197, d174, d185);
	xnor (d198, d171, d184);
	nor (d199, d155, d162);
	xor (d200, d171, d182);
	xnor (d201, d157, d169);
	xor (d202, d165, d178);
	buf (d203, d160);
	xnor (d204, d186);
	or (d205, d186, d188);
	or (d206, d155, d159);
	and (d207, d162, d181);
	not (d208, d107);
	buf (d209, d9);
	xor (d210, d158, d159);
	xor (d211, d171, d179);
	and (d212, d152, d173);
	xnor (d213, d160, d183);
	nor (d214, d157, d168);
	nand (d215, d171, d173);
	nor (d216, d161, d183);
	or (d217, d172, d187);
	xnor (d218, d170, d174);
	xor (d219, d155, d187);
	nand (d220, d152, d178);
	or (d221, d164, d169);
	buf (d222, d112);
	xnor (d223, d163, d185);
	or (d224, d166, d182);
	buf (d225, d21);
	nand (d226, d157, d170);
	and (d227, d157, d161);
	or (d228, d170, d188);
	not (d229, d147);
	xor (d230, d167, d180);
	xnor (d231, d154, d161);
	or (d232, d165, d179);
	or (d233, d165, d178);
	or (d234, d159, d162);
	and (d235, d168, d179);
	not (d236, d69);
	xor (d237, d191, d208);
	nand (d238, d201, d210);
	nor (d239, d218, d230);
	nand (d240, d196, d207);
	or (d241, d204, d208);
	xnor (d242, d213, d228);
	xor (d243, d200, d223);
	not (d244, d179);
	nor (d245, d198, d212);
	nor (d246, d189, d206);
	not (d247, d81);
	xor (d248, d228, d236);
	xnor (d249, d221, d227);
	nand (d250, d214, d231);
	xnor (d251, d191, d212);
	or (d252, d195, d208);
	buf (d253, d173);
	nor (d254, d194, d234);
	or (d255, d189, d202);
	xnor (d256, d198, d229);
	and (d257, d214, d226);
	xor (d258, d195, d223);
	xnor (d259, d196, d215);
	nor (d260, d194, d199);
	or (d261, d234, d235);
	not (d262, d224);
	not (d263, d138);
	xnor (d264, d201, d206);
	buf (d265, d135);
	xnor (d266, d201, d215);
	or (d267, d206, d231);
	buf (d268, d80);
	xor (d269, d189, d194);
	xor (d270, d203, d223);
	nand (d271, d216, d221);
	nand (d272, d196, d232);
	or (d273, d193, d196);
	nor (d274, d191, d208);
	or (d275, d205, d234);
	nand (d276, d193, d225);
	nand (d277, d224);
	or (d278, d191, d201);
	nor (d279, d200, d226);
	not (d280, d85);
	xor (d281, d203, d222);
	or (d282, d199, d219);
	and (d283, d198, d223);
	nor (d284, d256, d282);
	not (d285, d116);
	xnor (d286, d238, d280);
	nor (d287, d245, d250);
	nand (d288, d249, d254);
	nand (d289, d253, d272);
	buf (d290, d280);
	and (d291, d242, d279);
	nor (d292, d240, d252);
	xnor (d293, d238, d244);
	nor (d294, d237, d280);
	assign f1 = d287;
	assign f2 = d294;
	assign f3 = d285;
	assign f4 = d284;
	assign f5 = d284;
	assign f6 = d289;
	assign f7 = d289;
endmodule
