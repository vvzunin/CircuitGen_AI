module CCGRCG46( x0, x1, x2, f1, f2, f3, f4, f5, f6 );

	input x0, x1, x2;
	output f1, f2, f3, f4, f5, f6;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256;

	xor (d1, x0, x2);
	not (d2, x0);
	nand (d3, x1, x2);
	xor (d4, x1, x2);
	xnor (d5, x0, x1);
	not (d6, x1);
	nand (d7, x0, x2);
	xnor (d8, x1);
	and (d9, x0, x2);
	nor (d10, x1);
	or (d11, x2);
	and (d12, x1, x2);
	nand (d13, x2);
	buf (d14, x2);
	or (d15, x0);
	not (d16, x2);
	or (d17, x0, x2);
	nor (d18, x1, x2);
	xor (d19, x1);
	buf (d20, x0);
	xor (d21, x2);
	or (d22, x0, x2);
	or (d23, x0, x1);
	xor (d24, x0, x2);
	nand (d25, x1, x2);
	nor (d26, x0, x2);
	xnor (d27, x1, x2);
	xor (d28, x0, x1);
	nand (d29, x0, x2);
	xnor (d30, x0, x2);
	and (d31, x1);
	and (d32, x0, x1);
	xnor (d33, x0, x2);
	xnor (d34, x1, x2);
	buf (d35, x1);
	or (d36, x1, x2);
	nor (d37, x1, x2);
	nand (d38, x0, x1);
	nor (d39, x0, x2);
	and (d40, x0);
	xnor (d41, x0, x1);
	and (d42, x0, x1);
	and (d43, x1, x2);
	and (d44, d12, d32);
	buf (d45, d20);
	xor (d46, d18);
	nand (d47, d18, d39);
	nand (d48, d8, d33);
	buf (d49, d7);
	buf (d50, d3);
	buf (d51, d26);
	or (d52, d22, d33);
	xnor (d53, d6, d30);
	and (d54, d6, d41);
	nor (d55, d25, d32);
	not (d56, d15);
	nand (d57, d5, d14);
	buf (d58, d14);
	xnor (d59, d1, d41);
	not (d60, d22);
	nor (d61, d33, d41);
	nor (d62, d1, d9);
	or (d63, d9, d24);
	and (d64, d23, d31);
	or (d65, d19, d31);
	and (d66, d20, d29);
	not (d67, d23);
	xnor (d68, d11, d30);
	and (d69, d6, d28);
	xor (d70, d6, d13);
	nand (d71, d2, d38);
	nor (d72, d17);
	not (d73, d35);
	nand (d74, d20, d41);
	buf (d75, d12);
	xor (d76, d25, d28);
	xor (d77, d29, d36);
	and (d78, d33, d40);
	nor (d79, d6, d27);
	xor (d80, d37, d38);
	nand (d81, d27, d29);
	and (d82, d3, d24);
	xor (d83, d7, d43);
	xor (d84, d24, d34);
	and (d85, d26, d37);
	not (d86, d12);
	not (d87, d30);
	not (d88, d19);
	or (d89, d15, d33);
	xnor (d90, d9, d38);
	and (d91, d34, d36);
	xnor (d92, d17, d35);
	or (d93, d8, d36);
	nand (d94, d32, d38);
	and (d95, d3, d22);
	not (d96, d33);
	xor (d97, d69, d88);
	not (d98, d17);
	buf (d99, d37);
	buf (d100, d53);
	nand (d101, d54, d81);
	nand (d102, d97, d98);
	nand (d103, d98, d99);
	xnor (d104, d100, d101);
	nor (d105, d99, d100);
	not (d106, d31);
	not (d107, d48);
	or (d108, d97, d100);
	or (d109, d100, d101);
	xor (d110, d98, d100);
	nor (d111, d97, d101);
	xnor (d112, d99, d100);
	xor (d113, d98, d100);
	and (d114, d99);
	nand (d115, d98, d99);
	nor (d116, d97, d98);
	or (d117, d97, d98);
	nor (d118, d101);
	xor (d119, d97, d100);
	buf (d120, d82);
	buf (d121, d62);
	xnor (d122, d97, d99);
	and (d123, d99, d101);
	buf (d124, d51);
	and (d125, d98, d100);
	xor (d126, d101);
	and (d127, d100, d101);
	or (d128, d98);
	xor (d129, d98, d99);
	nor (d130, d99, d101);
	nand (d131, d97, d100);
	buf (d132, d87);
	xnor (d133, d99, d101);
	nand (d134, d97, d101);
	and (d135, d97, d98);
	buf (d136, d19);
	or (d137, d100);
	and (d138, d97, d100);
	nor (d139, d97, d100);
	or (d140, d98, d99);
	nor (d141, d98, d99);
	and (d142, d98, d101);
	xnor (d143, d97, d100);
	nand (d144, d100, d101);
	nor (d145, d98, d101);
	not (d146, d90);
	nand (d147, d98, d101);
	and (d148, d98, d99);
	xnor (d149, d97, d99);
	nand (d150, d99, d101);
	nand (d151, d97, d99);
	xor (d152, d99, d100);
	xor (d153, d99, d101);
	or (d154, d98, d99);
	or (d155, d98, d100);
	nor (d156, d98, d99);
	xnor (d157, d100);
	not (d158, d32);
	nor (d159, d100);
	and (d160, d97, d99);
	nor (d161, d97, d101);
	not (d162, d41);
	not (d163, d10);
	or (d164, d99, d101);
	nand (d165, d100, d101);
	or (d166, d97, d98);
	buf (d167, d49);
	xor (d168, d99, d100);
	xnor (d169, d98, d101);
	xor (d170, d100);
	buf (d171, d68);
	buf (d172, d57);
	nand (d173, d97, d101);
	and (d174, d141, d146);
	buf (d175, d97);
	not (d176, d120);
	nand (d177, d124, d146);
	buf (d178, d129);
	nor (d179, d136, d151);
	and (d180, d128, d149);
	xnor (d181, d107, d149);
	xnor (d182, d124, d130);
	xnor (d183, d122, d155);
	or (d184, d130, d137);
	not (d185, d55);
	nand (d186, d130, d141);
	nor (d187, d153, d172);
	xor (d188, d129, d162);
	xnor (d189, d115, d143);
	xnor (d190, d132, d149);
	nand (d191, d119, d155);
	and (d192, d119, d157);
	or (d193, d116, d162);
	xor (d194, d104, d157);
	not (d195, d93);
	xnor (d196, d161, d166);
	nand (d197, d141, d155);
	or (d198, d148, d167);
	nor (d199, d148, d154);
	xnor (d200, d103, d125);
	buf (d201, d79);
	xor (d202, d144, d156);
	and (d203, d103, d169);
	or (d204, d106, d170);
	nand (d205, d106, d146);
	and (d206, d156, d173);
	buf (d207, d132);
	xor (d208, d122, d172);
	xnor (d209, d124, d136);
	not (d210, d110);
	or (d211, d124, d163);
	xnor (d212, d108, d163);
	or (d213, d120, d168);
	nand (d214, d104, d149);
	xor (d215, d114, d140);
	or (d216, d144, d155);
	nor (d217, d113, d124);
	xor (d218, d134, d159);
	not (d219, d6);
	not (d220, d152);
	not (d221, d107);
	not (d222, d129);
	xnor (d223, d103, d112);
	not (d224, d126);
	xnor (d225, d102, d156);
	nand (d226, d139, d166);
	xnor (d227, d105, d170);
	nor (d228, d139, d172);
	or (d229, d107, d121);
	buf (d230, d84);
	not (d231, d165);
	nand (d232, d140, d147);
	or (d233, d154, d156);
	xnor (d234, d145, d153);
	not (d235, d28);
	nand (d236, d109, d139);
	nor (d237, d135, d144);
	not (d238, d128);
	nor (d239, d149, d157);
	and (d240, d111, d168);
	xnor (d241, d139, d141);
	not (d242, d100);
	buf (d243, d41);
	nor (d244, d116, d141);
	or (d245, d107, d137);
	xor (d246, d105, d172);
	and (d247, d134, d168);
	nor (d248, d128, d172);
	xnor (d249, d110, d152);
	xor (d250, d102, d154);
	not (d251, d61);
	not (d252, d139);
	xor (d253, d123, d151);
	xor (d254, d105, d125);
	xnor (d255, d153);
	nor (d256, d129);
	assign f1 = d237;
	assign f2 = d189;
	assign f3 = d206;
	assign f4 = d256;
	assign f5 = d187;
	assign f6 = d211;
endmodule
