module CCGRCG68( x0, x1, x2, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17 );

	input x0, x1, x2;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314, d315, d316;

	nor (d1, x0);
	and (d2, x0, x2);
	xor (d3, d1, d2);
	and (d4, d1, d2);
	nor (d5, d1, d2);
	or (d6, d1, d2);
	buf (d7, x0);
	nand (d8, d1, d2);
	xnor (d9, d2);
	buf (d10, d1);
	not (d11, x1);
	xnor (d12, d1, d2);
	or (d13, d1, d2);
	buf (d14, d2);
	xor (d15, d10, d11);
	xor (d16, d5, d7);
	xor (d17, d3);
	and (d18, d13, d14);
	or (d19, d6, d11);
	nor (d20, d4, d5);
	xnor (d21, d6, d9);
	and (d22, d12, d14);
	buf (d23, d11);
	not (d24, d5);
	nor (d25, d4);
	nor (d26, d9);
	not (d27, d1);
	buf (d28, d4);
	or (d29, d4, d10);
	or (d30, d11, d14);
	or (d31, d4, d12);
	xor (d32, d12, d13);
	xor (d33, d8, d13);
	xnor (d34, d4, d8);
	buf (d35, d8);
	and (d36, d3, d14);
	nand (d37, d11, d12);
	not (d38, d8);
	or (d39, d11, d14);
	not (d40, d13);
	xor (d41, d12, d14);
	and (d42, d4, d12);
	not (d43, d11);
	not (d44, d10);
	xor (d45, d3, d12);
	or (d46, d3, d5);
	not (d47, d4);
	or (d48, d3, d12);
	xnor (d49, d3, d7);
	buf (d50, d7);
	or (d51, d7, d12);
	nand (d52, d11, d13);
	nand (d53, d9, d14);
	nor (d54, d8, d13);
	and (d55, d7, d13);
	and (d56, d7, d13);
	or (d57, d8, d14);
	nor (d58, d3, d14);
	and (d59, d6, d9);
	or (d60, d3, d7);
	and (d61, d3, d9);
	and (d62, d3, d5);
	or (d63, d10, d14);
	xor (d64, d12, d14);
	xor (d65, d6, d10);
	and (d66, d10, d12);
	nor (d67, d7, d10);
	and (d68, d5, d8);
	nand (d69, d7, d14);
	and (d70, d4, d9);
	xor (d71, d3, d6);
	not (d72, d6);
	and (d73, d4, d14);
	nand (d74, d10, d13);
	nor (d75, d8, d14);
	nand (d76, d5, d9);
	nor (d77, d6, d14);
	nand (d78, d7, d10);
	or (d79, d12);
	buf (d80, d14);
	and (d81, d4, d12);
	or (d82, d5, d13);
	nand (d83, d8, d14);
	or (d84, d5, d14);
	nand (d85, d4, d7);
	nor (d86, d6, d7);
	nor (d87, d9, d13);
	nor (d88, d8, d10);
	xnor (d89, d5, d7);
	nor (d90, d4, d8);
	nor (d91, d6, d10);
	xnor (d92, d4, d12);
	xor (d93, d6, d12);
	and (d94, d9, d11);
	and (d95, d3, d10);
	nand (d96, d3, d13);
	xnor (d97, d27, d77);
	nand (d98, d51, d90);
	xnor (d99, d23, d72);
	xor (d100, d36, d66);
	or (d101, d23, d58);
	or (d102, d41, d82);
	and (d103, d31, d83);
	xor (d104, d31, d60);
	nor (d105, d87, d91);
	nor (d106, d32, d59);
	not (d107, d36);
	xnor (d108, d31, d69);
	buf (d109, d76);
	buf (d110, d91);
	buf (d111, d26);
	or (d112, d58, d59);
	and (d113, d55, d76);
	not (d114, d75);
	xnor (d115, d98, d112);
	not (d116, d48);
	not (d117, d110);
	buf (d118, d87);
	xnor (d119, d107, d113);
	nor (d120, d105, d108);
	and (d121, d101, d106);
	and (d122, d101, d104);
	buf (d123, d37);
	nor (d124, d105, d107);
	not (d125, d68);
	nor (d126, d106, d113);
	buf (d127, d68);
	nor (d128, d104, d112);
	buf (d129, d23);
	xnor (d130, d105);
	xnor (d131, d101, d103);
	nor (d132, d98, d106);
	buf (d133, d22);
	or (d134, d100, d113);
	buf (d135, d110);
	buf (d136, d65);
	xor (d137, d114, d126);
	xor (d138, d124, d126);
	and (d139, d120, d121);
	buf (d140, d132);
	nand (d141, d126, d129);
	and (d142, d115, d116);
	buf (d143, d92);
	xor (d144, d125, d128);
	not (d145, d128);
	and (d146, d125, d130);
	buf (d147, d15);
	xnor (d148, d117, d132);
	buf (d149, d129);
	nand (d150, d125, d132);
	xnor (d151, d118, d134);
	and (d152, d119, d131);
	xor (d153, d114, d121);
	or (d154, d119, d124);
	xnor (d155, d124, d126);
	or (d156, d116, d134);
	not (d157, d86);
	nand (d158, d118, d133);
	not (d159, d38);
	buf (d160, d100);
	xor (d161, d127, d134);
	or (d162, d123, d131);
	xor (d163, d119, d128);
	xnor (d164, d114, d124);
	or (d165, d119, d123);
	and (d166, d128, d133);
	nor (d167, d123, d131);
	xor (d168, d120, d125);
	and (d169, d127, d134);
	xnor (d170, d115);
	and (d171, d119, d122);
	xnor (d172, d117, d127);
	or (d173, d128, d129);
	xor (d174, d123, d131);
	xor (d175, d122, d129);
	nand (d176, d119, d122);
	nor (d177, d114, d116);
	nand (d178, d119, d132);
	or (d179, d118, d124);
	buf (d180, d52);
	nor (d181, d115, d130);
	and (d182, d120, d129);
	nand (d183, d124, d125);
	or (d184, d120, d125);
	xor (d185, d116, d131);
	nand (d186, d118, d119);
	not (d187, d115);
	nand (d188, d127, d131);
	buf (d189, d78);
	not (d190, d120);
	xor (d191, d118, d124);
	not (d192, d112);
	not (d193, d52);
	xnor (d194, d123, d127);
	xnor (d195, d123, d131);
	xor (d196, d122, d126);
	xor (d197, d120, d125);
	not (d198, d113);
	not (d199, d108);
	nand (d200, d114, d115);
	not (d201, d77);
	not (d202, d17);
	or (d203, d128, d129);
	and (d204, d114, d133);
	not (d205, d57);
	xor (d206, d118, d127);
	nor (d207, d115, d125);
	and (d208, d116, d119);
	nor (d209, d115, d117);
	nor (d210, d123, d127);
	or (d211, d118, d125);
	nand (d212, d116, d127);
	and (d213, d120, d133);
	nand (d214, d121, d126);
	buf (d215, d34);
	buf (d216, d206);
	not (d217, d114);
	and (d218, d158, d169);
	buf (d219, d176);
	nand (d220, d181, d184);
	xor (d221, d182, d207);
	or (d222, d184, d204);
	and (d223, d148, d192);
	nor (d224, d165, d171);
	buf (d225, d130);
	and (d226, d149, d166);
	xnor (d227, d179, d194);
	and (d228, d175, d176);
	and (d229, d168, d214);
	and (d230, d157, d201);
	buf (d231, d173);
	or (d232, d156, d211);
	and (d233, d156, d168);
	xor (d234, d156, d162);
	not (d235, d98);
	or (d236, d155, d207);
	nand (d237, d135, d161);
	nand (d238, d185, d199);
	or (d239, d186, d197);
	xor (d240, d163, d211);
	or (d241, d191, d197);
	xnor (d242, d141, d176);
	nand (d243, d144, d213);
	xor (d244, d167, d170);
	or (d245, d141, d192);
	xnor (d246, d136, d183);
	and (d247, d207, d211);
	not (d248, d178);
	xnor (d249, d221, d229);
	and (d250, d234, d240);
	xnor (d251, d220, d224);
	or (d252, d231, d243);
	nor (d253, d233, d246);
	buf (d254, d10);
	and (d255, d219, d246);
	or (d256, d219, d245);
	nand (d257, d236, d239);
	or (d258, d233, d246);
	xnor (d259, d243, d245);
	or (d260, d225, d231);
	xnor (d261, d232, d238);
	or (d262, d232, d246);
	nand (d263, d238, d245);
	xor (d264, d227, d242);
	and (d265, d233, d243);
	nor (d266, d226, d233);
	nand (d267, d222, d228);
	buf (d268, d75);
	xor (d269, d222, d247);
	nor (d270, d216, d218);
	nand (d271, d227, d241);
	buf (d272, d111);
	buf (d273, d140);
	xor (d274, d228, d241);
	or (d275, d221, d230);
	and (d276, d259, d273);
	not (d277, d19);
	nand (d278, d253, d270);
	xor (d279, d262, d268);
	xnor (d280, d259, d264);
	xor (d281, d251, d260);
	nor (d282, d264, d270);
	nand (d283, d266, d270);
	and (d284, d268, d269);
	nor (d285, d265, d271);
	xor (d286, d259, d275);
	nand (d287, d256, d270);
	buf (d288, d156);
	not (d289, d135);
	xor (d290, d255);
	and (d291, d252, d274);
	buf (d292, d146);
	xor (d293, d254, d274);
	xnor (d294, d265, d272);
	xor (d295, d253, d261);
	nand (d296, d271);
	and (d297, d265, d266);
	buf (d298, d193);
	buf (d299, d205);
	nor (d300, d252, d254);
	not (d301, d129);
	nand (d302, d259, d261);
	buf (d303, d40);
	not (d304, d84);
	xnor (d305, d270, d273);
	xnor (d306, d260, d262);
	and (d307, d260, d264);
	or (d308, d262, d274);
	nand (d309, d256, d265);
	nor (d310, d256, d260);
	xnor (d311, d267, d275);
	nand (d312, d253, d270);
	xor (d313, d256, d263);
	nor (d314, d250, d271);
	or (d315, d267);
	or (d316, d252, d275);
	assign f1 = d311;
	assign f2 = d277;
	assign f3 = d310;
	assign f4 = d306;
	assign f5 = d286;
	assign f6 = d290;
	assign f7 = d292;
	assign f8 = d308;
	assign f9 = d289;
	assign f10 = d279;
	assign f11 = d278;
	assign f12 = d277;
	assign f13 = d284;
	assign f14 = d315;
	assign f15 = d290;
	assign f16 = d293;
	assign f17 = d282;
endmodule
