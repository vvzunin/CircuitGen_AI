module CCGRCG58( x0, x1, x2, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12 );

	input x0, x1, x2;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314, d315, d316, d317, d318, d319, d320, d321, d322, d323, d324, d325, d326, d327, d328, d329, d330, d331, d332, d333, d334, d335, d336, d337, d338, d339, d340, d341, d342, d343, d344, d345, d346, d347, d348, d349, d350, d351, d352, d353, d354, d355, d356, d357, d358, d359, d360, d361, d362, d363, d364, d365, d366;

	or (d1, x0, x2);
	not (d2, x2);
	and (d3, x2);
	nand (d4, x0);
	or (d5, x1, x2);
	nor (d6, x1, x2);
	xnor (d7, x0, x1);
	nand (d8, x0, x1);
	and (d9, x0, x1);
	nor (d10, x0, x2);
	and (d11, x0, x2);
	buf (d12, x2);
	xnor (d13, x0);
	xnor (d14, x0, x2);
	xor (d15, x0, x1);
	buf (d16, x1);
	not (d17, x1);
	xnor (d18, x0, x2);
	xor (d19, x1, x2);
	or (d20, x1, x2);
	nor (d21, x1, x2);
	buf (d22, x0);
	or (d23, x0, x2);
	and (d24, d8, d9);
	and (d25, d1, d7);
	buf (d26, d15);
	buf (d27, d7);
	xor (d28, d1, d20);
	xor (d29, d17, d23);
	nand (d30, d6, d21);
	xor (d31, d7, d18);
	nand (d32, d1, d15);
	xnor (d33, d12, d15);
	not (d34, d13);
	xnor (d35, d9, d13);
	not (d36, d19);
	or (d37, d3, d5);
	nor (d38, d2, d18);
	not (d39, d1);
	and (d40, d2, d5);
	buf (d41, d19);
	or (d42, d11, d13);
	nor (d43, d11, d23);
	nor (d44, d2, d4);
	and (d45, d5, d16);
	buf (d46, d16);
	xor (d47, d1, d7);
	not (d48, d2);
	nor (d49, d18, d23);
	nand (d50, d4, d5);
	and (d51, d18, d21);
	nor (d52, d14, d18);
	nor (d53, d1, d4);
	not (d54, x0);
	xor (d55, d9);
	nor (d56, d3, d6);
	or (d57, d10, d19);
	buf (d58, d5);
	nor (d59, d23);
	xnor (d60, d1);
	not (d61, d15);
	or (d62, d11, d16);
	nand (d63, d8, d14);
	nand (d64, d9, d23);
	nand (d65, d12, d17);
	not (d66, d22);
	or (d67, d9, d14);
	not (d68, d8);
	nor (d69, d8, d15);
	not (d70, d12);
	xor (d71, d5, d9);
	buf (d72, d18);
	nand (d73, d10, d17);
	or (d74, d1, d12);
	nand (d75, d1, d12);
	and (d76, d9, d20);
	nor (d77, d2, d21);
	not (d78, d9);
	not (d79, d10);
	nand (d80, d2, d3);
	buf (d81, d13);
	xnor (d82, d68, d73);
	and (d83, d31, d33);
	nor (d84, d40, d73);
	xor (d85, d52, d54);
	or (d86, d36, d65);
	buf (d87, d6);
	and (d88, d32, d37);
	and (d89, d56, d65);
	xor (d90, d50, d58);
	nand (d91, d33, d57);
	xor (d92, d56, d78);
	nand (d93, d40, d77);
	xnor (d94, d32, d33);
	xor (d95, d32, d62);
	xnor (d96, d42, d71);
	or (d97, d85, d96);
	not (d98, d54);
	not (d99, d73);
	nor (d100, d84, d94);
	nor (d101, d92, d94);
	buf (d102, d93);
	nor (d103, d84, d92);
	buf (d104, d31);
	nand (d105, d86, d87);
	nand (d106, d90, d92);
	xor (d107, d81, d95);
	xor (d108, d85, d89);
	xnor (d109, d89, d90);
	nor (d110, d85, d87);
	xor (d111, d91, d95);
	xnor (d112, d83, d85);
	nor (d113, d85, d86);
	nor (d114, d83, d86);
	xnor (d115, d89, d90);
	or (d116, d83, d94);
	xnor (d117, d103, d114);
	not (d118, d84);
	or (d119, d107, d111);
	nor (d120, d112, d114);
	nand (d121, d105, d107);
	nor (d122, d108, d109);
	xor (d123, d107, d115);
	not (d124, d27);
	and (d125, d103, d113);
	xnor (d126, d109, d113);
	nor (d127, d100, d108);
	xnor (d128, d114, d116);
	and (d129, d105);
	not (d130, d80);
	buf (d131, d20);
	xnor (d132, d114);
	nand (d133, d98, d109);
	nand (d134, d100, d103);
	nand (d135, d111, d114);
	xor (d136, d99, d105);
	or (d137, d110, d111);
	xor (d138, d113);
	buf (d139, d10);
	xor (d140, d105, d110);
	nor (d141, d100, d112);
	nor (d142, d98, d111);
	nor (d143, d131, d138);
	nand (d144, d123, d141);
	xor (d145, d122, d133);
	not (d146, d106);
	nor (d147, d125, d126);
	xor (d148, d121, d131);
	xor (d149, d137, d140);
	or (d150, d117, d134);
	not (d151, d112);
	or (d152, d138, d141);
	nand (d153, d119, d138);
	nand (d154, d123, d134);
	xor (d155, d118, d119);
	and (d156, d124, d140);
	and (d157, d129, d139);
	and (d158, d133, d139);
	xor (d159, d123, d138);
	nand (d160, d126, d129);
	not (d161, d135);
	not (d162, d77);
	or (d163, d129, d133);
	not (d164, d64);
	xor (d165, d124, d138);
	or (d166, d125, d127);
	nor (d167, d123, d126);
	nor (d168, d119, d127);
	or (d169, d118, d126);
	or (d170, d137, d141);
	xnor (d171, d118, d128);
	xor (d172, d132, d137);
	not (d173, d31);
	xnor (d174, d132);
	buf (d175, d134);
	xor (d176, d128, d141);
	or (d177, d118, d127);
	nor (d178, d134, d140);
	not (d179, d103);
	and (d180, d123, d133);
	xor (d181, d133, d134);
	xor (d182, d138, d139);
	xor (d183, d133, d134);
	nor (d184, d132, d141);
	buf (d185, d102);
	nand (d186, d121, d140);
	nand (d187, d122, d127);
	buf (d188, d133);
	xor (d189, d120, d122);
	xor (d190, d119, d141);
	or (d191, d130, d134);
	xor (d192, d123, d131);
	xor (d193, d130, d137);
	and (d194, d118, d130);
	nand (d195, d140);
	xnor (d196, d120, d137);
	nand (d197, d123, d132);
	and (d198, d120, d129);
	xor (d199, d121, d123);
	xor (d200, d127, d142);
	or (d201, d117, d136);
	and (d202, d154, d163);
	nor (d203, d165, d168);
	xor (d204, d173, d183);
	nand (d205, d149, d167);
	nor (d206, d201);
	buf (d207, d195);
	not (d208, d93);
	buf (d209, d14);
	or (d210, d150, d194);
	not (d211, d167);
	and (d212, d146, d161);
	nand (d213, d147, d176);
	or (d214, d143, d174);
	and (d215, d162, d180);
	nand (d216, d181, d188);
	xnor (d217, d160, d171);
	nand (d218, d147, d171);
	nor (d219, d165, d185);
	nor (d220, d155, d191);
	buf (d221, d175);
	or (d222, d167, d183);
	nand (d223, d173, d191);
	or (d224, d165, d174);
	xnor (d225, d176, d187);
	buf (d226, d48);
	xor (d227, d185, d198);
	nand (d228, d153, d183);
	not (d229, d78);
	nand (d230, d161, d197);
	and (d231, d176, d190);
	not (d232, d88);
	xnor (d233, d157, d160);
	xnor (d234, d185, d186);
	nand (d235, d164, d176);
	nand (d236, d167, d175);
	xnor (d237, d146, d186);
	not (d238, d142);
	not (d239, d82);
	nor (d240, d155, d178);
	and (d241, d192, d198);
	and (d242, d192, d197);
	and (d243, d152, d179);
	and (d244, d187, d196);
	nor (d245, d186, d192);
	buf (d246, d183);
	xnor (d247, d193, d201);
	xnor (d248, d156, d190);
	nor (d249, d145, d171);
	and (d250, d164, d169);
	xor (d251, d147, d170);
	nor (d252, d184, d187);
	or (d253, d172, d196);
	xnor (d254, d182, d189);
	not (d255, d158);
	not (d256, d72);
	buf (d257, d72);
	or (d258, d159, d190);
	or (d259, d193, d195);
	xor (d260, d162, d183);
	not (d261, d134);
	xor (d262, d147, d185);
	not (d263, d173);
	xnor (d264, d152, d194);
	xnor (d265, d164, d168);
	xnor (d266, d167, d191);
	or (d267, d161, d162);
	nand (d268, d162, d178);
	xnor (d269, d165, d187);
	xor (d270, d193, d198);
	buf (d271, d141);
	not (d272, d75);
	not (d273, d42);
	and (d274, d151, d193);
	not (d275, d190);
	xnor (d276, d170, d172);
	and (d277, d157, d168);
	buf (d278, d90);
	xnor (d279, d150, d191);
	and (d280, d220, d223);
	nor (d281, d203, d271);
	and (d282, d224);
	buf (d283, d240);
	not (d284, d258);
	xor (d285, d259, d262);
	not (d286, d206);
	or (d287, d209, d212);
	not (d288, d6);
	and (d289, d209, d230);
	xnor (d290, d257, d269);
	xor (d291, d242, d265);
	xor (d292, d204, d236);
	not (d293, d176);
	and (d294, d260, d274);
	xor (d295, d251, d274);
	xnor (d296, d227, d265);
	or (d297, d207, d224);
	xor (d298, d258, d261);
	not (d299, d138);
	xnor (d300, d255, d266);
	xnor (d301, d225, d277);
	not (d302, d223);
	nor (d303, d219, d262);
	nand (d304, d211, d267);
	and (d305, d224, d247);
	xnor (d306, d241, d270);
	and (d307, d204, d249);
	nor (d308, d212, d225);
	not (d309, d210);
	and (d310, d235, d272);
	xnor (d311, d249, d275);
	buf (d312, d273);
	not (d313, d217);
	xnor (d314, d223, d250);
	nor (d315, d207, d279);
	nor (d316, d217, d278);
	not (d317, d18);
	or (d318, d233, d244);
	xnor (d319, d276, d277);
	not (d320, d4);
	nor (d321, d297, d318);
	xor (d322, d282, d308);
	or (d323, d282, d292);
	xnor (d324, d286, d291);
	buf (d325, d264);
	xnor (d326, d283, d300);
	not (d327, d171);
	xor (d328, d287, d300);
	xor (d329, d298, d306);
	xnor (d330, d304, d316);
	buf (d331, d181);
	and (d332, d286, d314);
	and (d333, d285, d307);
	nand (d334, d285, d308);
	not (d335, d123);
	xor (d336, d299, d310);
	nand (d337, d304, d310);
	or (d338, d289, d296);
	xor (d339, d295, d296);
	or (d340, d286, d311);
	or (d341, d282, d293);
	buf (d342, d276);
	nand (d343, d281, d316);
	xnor (d344, d280, d316);
	or (d345, d297, d319);
	xor (d346, d314, d316);
	nor (d347, d280, d297);
	or (d348, d302, d319);
	buf (d349, d224);
	xor (d350, d309);
	nand (d351, d302);
	xor (d352, d312, d317);
	xor (d353, d315, d318);
	xor (d354, d291, d304);
	xnor (d355, d304, d305);
	nand (d356, d282, d315);
	nor (d357, d288, d309);
	nor (d358, d296, d312);
	not (d359, d219);
	or (d360, d284, d306);
	xor (d361, d282, d284);
	nand (d362, d306, d313);
	buf (d363, d194);
	or (d364, d288, d291);
	xnor (d365, d292, d304);
	and (d366, d307, d317);
	assign f1 = d325;
	assign f2 = d334;
	assign f3 = d325;
	assign f4 = d345;
	assign f5 = d322;
	assign f6 = d320;
	assign f7 = d325;
	assign f8 = d366;
	assign f9 = d322;
	assign f10 = d346;
	assign f11 = d331;
	assign f12 = d348;
endmodule
