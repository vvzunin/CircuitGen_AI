module CCGRCG141( x0, x1, x2, x3, x4, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15 );

	input x0, x1, x2, x3, x4;
	output f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15;

	wire d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314, d315, d316, d317, d318, d319, d320, d321, d322, d323, d324, d325, d326, d327, d328, d329, d330, d331, d332, d333, d334, d335, d336, d337, d338, d339, d340, d341, d342, d343, d344, d345, d346, d347, d348, d349, d350, d351, d352, d353, d354, d355, d356, d357, d358, d359, d360, d361, d362, d363, d364, d365, d366, d367, d368, d369, d370, d371, d372, d373, d374, d375, d376, d377, d378, d379, d380, d381, d382, d383, d384, d385, d386, d387, d388, d389, d390, d391, d392, d393, d394, d395, d396, d397, d398, d399, d400, d401, d402, d403, d404, d405, d406, d407, d408, d409, d410, d411, d412, d413, d414, d415, d416, d417, d418, d419, d420, d421, d422, d423, d424, d425, d426, d427, d428, d429, d430, d431, d432, d433, d434, d435, d436, d437, d438, d439, d440, d441, d442, d443, d444, d445, d446, d447, d448, d449, d450, d451, d452, d453, d454, d455, d456, d457, d458, d459, d460, d461, d462, d463, d464, d465, d466, d467, d468, d469, d470, d471, d472, d473, d474, d475, d476, d477, d478, d479, d480, d481, d482, d483, d484, d485, d486, d487, d488, d489, d490, d491, d492, d493, d494, d495, d496, d497, d498, d499, d500, d501, d502, d503, d504, d505, d506, d507, d508, d509, d510, d511, d512, d513, d514, d515, d516, d517, d518;

	nand (d1, x1, x2);
	buf (d2, x4);
	xor (d3, x2, x3);
	or (d4, x1, x4);
	buf (d5, x2);
	or (d6, x3, x4);
	buf (d7, x0);
	or (d8, x2, x4);
	or (d9, x1, x2);
	not (d10, x2);
	and (d11, x0, x3);
	not (d12, x3);
	or (d13, x1, x3);
	nor (d14, x3, x4);
	or (d15, x3);
	xnor (d16, x1);
	or (d17, x0, x4);
	nor (d18, x2, x3);
	xnor (d19, x2);
	xor (d20, x1, x4);
	xor (d21, x1, x4);
	nand (d22, x3, x4);
	and (d23, x0, x1);
	not (d24, x4);
	xnor (d25, x0, x2);
	and (d26, x3);
	nand (d27, x2, x3);
	nor (d28, x0);
	nor (d29, x4);
	xor (d30, x1);
	xnor (d31, x3);
	not (d32, x1);
	nor (d33, x1, x2);
	xnor (d34, x1, x2);
	nand (d35, x1, x4);
	or (d36, x0);
	and (d37, x1);
	xnor (d38, x0, x3);
	xnor (d39, x0);
	and (d40, x0, x1);
	and (d41, x4);
	nand (d42, x1, x2);
	nand (d43, x0, x3);
	buf (d44, x3);
	nor (d45, x2, x4);
	and (d46, x2, x4);
	not (d47, x0);
	or (d48, x4);
	and (d49, x2, x3);
	or (d50, d13, d30);
	and (d51, d2, d6);
	nand (d52, d5, d13);
	not (d53, d25);
	xnor (d54, d1, d17);
	not (d55, d36);
	nand (d56, d5, d28);
	xnor (d57, d27, d49);
	nand (d58, d54, d56);
	or (d59, d56, d57);
	nor (d60, d50, d56);
	nor (d61, d56);
	xor (d62, d51);
	or (d63, d51);
	nor (d64, d54, d57);
	nor (d65, d55, d56);
	not (d66, d32);
	nor (d67, d50, d52);
	or (d68, d54, d55);
	and (d69, d50, d55);
	xor (d70, d51, d56);
	or (d71, d54);
	xor (d72, d50, d53);
	nand (d73, d54, d56);
	and (d74, d51, d57);
	xnor (d75, d52, d54);
	xor (d76, d52, d57);
	buf (d77, d5);
	buf (d78, d31);
	buf (d79, d45);
	xor (d80, d50, d52);
	nor (d81, d50, d54);
	nand (d82, d50, d57);
	or (d83, d50, d51);
	and (d84, d50, d52);
	buf (d85, d14);
	and (d86, d50, d57);
	nand (d87, d50, d56);
	xnor (d88, d50, d53);
	or (d89, d52, d56);
	or (d90, d50, d53);
	and (d91, d52, d57);
	not (d92, d42);
	xnor (d93, d53, d57);
	nand (d94, d52);
	and (d95, d54, d56);
	nand (d96, d54);
	xnor (d97, d51, d54);
	xor (d98, d55, d56);
	xor (d99, d52, d55);
	and (d100, d50, d57);
	not (d101, d38);
	nor (d102, d52, d54);
	not (d103, d26);
	xnor (d104, d53, d54);
	nand (d105, d51, d56);
	buf (d106, d3);
	buf (d107, d54);
	and (d108, d52, d53);
	and (d109, d52, d54);
	or (d110, d51, d52);
	xnor (d111, d51, d56);
	xor (d112, d50, d54);
	nor (d113, d51, d55);
	xor (d114, d53);
	nor (d115, d54);
	nor (d116, d54, d57);
	nand (d117, d51, d56);
	xor (d118, d53, d55);
	not (d119, d12);
	nand (d120, d51, d52);
	xor (d121, d55);
	nand (d122, d50);
	nor (d123, d59, d84);
	xor (d124, d109, d117);
	buf (d125, d115);
	and (d126, d78, d120);
	xnor (d127, d76, d100);
	xnor (d128, d73, d84);
	xnor (d129, d83, d99);
	xor (d130, d69, d108);
	xnor (d131, d73, d122);
	xor (d132, d72, d90);
	xnor (d133, d95, d108);
	nor (d134, d93, d119);
	nand (d135, d73, d104);
	xor (d136, d62, d118);
	nor (d137, d59, d68);
	xor (d138, d82, d118);
	not (d139, d11);
	or (d140, d92, d115);
	nand (d141, d63, d117);
	nor (d142, d105, d114);
	and (d143, d74, d98);
	nand (d144, d62, d120);
	buf (d145, d122);
	nor (d146, d59, d97);
	and (d147, d80, d93);
	buf (d148, d83);
	nor (d149, d79, d84);
	buf (d150, d23);
	nand (d151, d83, d121);
	nor (d152, d101, d116);
	or (d153, d72, d94);
	nor (d154, d102, d122);
	nor (d155, d143, d152);
	xnor (d156, d123, d146);
	buf (d157, d152);
	xnor (d158, d131, d132);
	and (d159, d149, d154);
	and (d160, d134, d143);
	xnor (d161, d125, d137);
	not (d162, d18);
	buf (d163, d12);
	or (d164, d124, d137);
	xor (d165, d124, d134);
	nor (d166, d139, d148);
	or (d167, d126, d129);
	or (d168, d133, d134);
	nand (d169, d130, d142);
	not (d170, d130);
	and (d171, d123, d153);
	xor (d172, d147, d149);
	nand (d173, d126, d149);
	not (d174, d7);
	buf (d175, d105);
	and (d176, d126, d147);
	or (d177, d130, d141);
	not (d178, d34);
	nand (d179, d130, d137);
	not (d180, d58);
	xnor (d181, d140, d153);
	buf (d182, d106);
	nor (d183, d142, d152);
	xor (d184, d141, d145);
	or (d185, d131, d140);
	nand (d186, d125, d145);
	not (d187, d148);
	nand (d188, d125, d132);
	nand (d189, d156, d169);
	not (d190, d40);
	and (d191, d159, d162);
	and (d192, d171, d174);
	buf (d193, d44);
	xor (d194, d169, d173);
	xnor (d195, d168, d171);
	xor (d196, d175, d182);
	nand (d197, d174, d176);
	buf (d198, d51);
	not (d199, d52);
	nand (d200, d173, d178);
	buf (d201, d90);
	nor (d202, d158, d163);
	or (d203, d159, d161);
	or (d204, d158, d160);
	nor (d205, d172, d174);
	xnor (d206, d166, d170);
	buf (d207, d10);
	or (d208, d177, d179);
	buf (d209, d102);
	xor (d210, d165, d169);
	and (d211, d161, d168);
	nor (d212, d157, d176);
	not (d213, d24);
	xor (d214, d173, d184);
	or (d215, d186, d188);
	not (d216, d19);
	and (d217, d178, d188);
	not (d218, d110);
	xnor (d219, d157, d178);
	nand (d220, d162, d172);
	xor (d221, d157, d177);
	or (d222, d158, d175);
	or (d223, d160, d173);
	buf (d224, d184);
	and (d225, d163, d175);
	nor (d226, d158, d186);
	not (d227, d169);
	xor (d228, d166, d187);
	buf (d229, d163);
	buf (d230, d145);
	xnor (d231, d160, d161);
	buf (d232, d142);
	and (d233, d158, d163);
	nand (d234, d155, d182);
	xnor (d235, d161, d187);
	xnor (d236, d175, d182);
	xor (d237, d174, d180);
	buf (d238, d171);
	buf (d239, d64);
	xor (d240, d155, d167);
	not (d241, d188);
	xor (d242, d163, d168);
	nor (d243, d165, d181);
	not (d244, d86);
	xnor (d245, d158, d161);
	nor (d246, d174, d181);
	not (d247, d77);
	xnor (d248, d159, d176);
	or (d249, d155, d170);
	nor (d250, d158, d160);
	or (d251, d160, d163);
	xnor (d252, d168, d180);
	xor (d253, d160, d172);
	not (d254, d93);
	or (d255, d170, d180);
	buf (d256, d25);
	buf (d257, d41);
	nand (d258, d184, d188);
	and (d259, d181, d187);
	buf (d260, d40);
	or (d261, d162, d186);
	nor (d262, d172, d173);
	nor (d263, d155, d177);
	nand (d264, d159, d167);
	nand (d265, d158, d179);
	xnor (d266, d173, d187);
	nand (d267, d170, d177);
	xor (d268, d179, d183);
	not (d269, d129);
	not (d270, d81);
	or (d271, d172, d181);
	and (d272, d164, d176);
	xnor (d273, d168, d181);
	xor (d274, d172, d173);
	and (d275, d163, d180);
	not (d276, d158);
	and (d277, d158, d168);
	nand (d278, d155, d156);
	or (d279, d157, d158);
	not (d280, d75);
	xnor (d281, d218, d223);
	nor (d282, d226, d259);
	buf (d283, d158);
	nor (d284, d260, d279);
	and (d285, d192, d227);
	not (d286, d10);
	nor (d287, d192, d217);
	xor (d288, d248, d261);
	xnor (d289, d223, d260);
	xor (d290, d231, d258);
	and (d291, d199, d206);
	nand (d292, d194, d199);
	and (d293, d195, d254);
	xor (d294, d257, d271);
	and (d295, d194, d215);
	xor (d296, d224, d231);
	nor (d297, d199, d265);
	and (d298, d216, d245);
	xnor (d299, d231, d263);
	and (d300, d193, d254);
	not (d301, d233);
	not (d302, d159);
	and (d303, d202, d253);
	and (d304, d233, d260);
	nor (d305, d247, d276);
	or (d306, d230, d236);
	xor (d307, d201, d220);
	xnor (d308, d206, d244);
	xor (d309, d225, d269);
	nor (d310, d249, d261);
	not (d311, d98);
	xor (d312, d235, d260);
	nor (d313, d192, d231);
	or (d314, d247, d262);
	nor (d315, d210, d255);
	nand (d316, d257, d272);
	nor (d317, d205, d217);
	or (d318, d274, d279);
	buf (d319, d252);
	nor (d320, d264, d276);
	or (d321, d193, d256);
	xnor (d322, d207, d248);
	nand (d323, d258, d277);
	xnor (d324, d191, d277);
	nor (d325, d210, d233);
	xnor (d326, d253, d259);
	not (d327, d92);
	and (d328, d209, d274);
	xnor (d329, d197, d267);
	nor (d330, d198, d237);
	xor (d331, d199, d253);
	nand (d332, d295, d330);
	buf (d333, d131);
	xnor (d334, d286, d311);
	xnor (d335, d304, d330);
	xnor (d336, d280, d311);
	not (d337, d164);
	xor (d338, d299, d310);
	xnor (d339, d284, d323);
	not (d340, d227);
	or (d341, d281, d326);
	or (d342, d312, d331);
	and (d343, d282, d299);
	xnor (d344, d296, d302);
	xor (d345, d288, d298);
	nor (d346, d283, d305);
	nand (d347, d310, d320);
	or (d348, d290, d319);
	nand (d349, d312, d320);
	and (d350, d284, d305);
	nand (d351, d292, d307);
	xor (d352, d302, d311);
	not (d353, d207);
	nand (d354, d290, d307);
	buf (d355, d237);
	nand (d356, d284, d328);
	nor (d357, d315, d319);
	and (d358, d293, d295);
	nor (d359, d284, d331);
	xor (d360, d280, d285);
	nor (d361, d324, d330);
	nand (d362, d286, d326);
	xnor (d363, d309, d313);
	xor (d364, d311, d322);
	xor (d365, d308, d316);
	nand (d366, d302, d324);
	buf (d367, d214);
	not (d368, d206);
	nand (d369, d292, d293);
	xor (d370, d286, d305);
	and (d371, d286, d330);
	not (d372, d142);
	xnor (d373, d294, d309);
	nor (d374, d284, d287);
	xor (d375, d297, d324);
	xor (d376, d284, d313);
	or (d377, d301, d309);
	and (d378, d282, d323);
	xnor (d379, d294, d305);
	and (d380, d319, d324);
	buf (d381, d34);
	buf (d382, d310);
	buf (d383, d177);
	or (d384, d293, d305);
	xor (d385, d296, d317);
	xnor (d386, d288, d296);
	not (d387, d187);
	xor (d388, d384, d386);
	buf (d389, d69);
	nor (d390, d354, d365);
	xnor (d391, d370, d381);
	xor (d392, d355, d369);
	or (d393, d356, d374);
	and (d394, d347, d377);
	nor (d395, d377, d379);
	xnor (d396, d335, d364);
	or (d397, d353, d356);
	nor (d398, d355, d368);
	or (d399, d347, d380);
	or (d400, d349, d355);
	xnor (d401, d354, d384);
	buf (d402, d73);
	nor (d403, d334, d368);
	nand (d404, d340, d368);
	xor (d405, d376, d377);
	xnor (d406, d343, d350);
	buf (d407, d215);
	and (d408, d337, d372);
	xor (d409, d350, d369);
	nand (d410, d344, d351);
	nor (d411, d340, d361);
	not (d412, d14);
	xor (d413, d347, d352);
	and (d414, d349, d379);
	or (d415, d354, d380);
	xor (d416, d337, d362);
	nand (d417, d349, d371);
	xor (d418, d365, d384);
	xnor (d419, d341, d350);
	and (d420, d350, d382);
	xor (d421, d342, d374);
	xnor (d422, d379, d380);
	not (d423, d369);
	buf (d424, d343);
	nand (d425, d361, d362);
	buf (d426, d239);
	xor (d427, d349, d352);
	not (d428, d141);
	xor (d429, d357, d379);
	and (d430, d352, d358);
	nor (d431, d360, d373);
	or (d432, d369, d370);
	and (d433, d384, d387);
	nor (d434, d366, d368);
	nand (d435, d359, d370);
	nand (d436, d336, d347);
	xnor (d437, d355, d367);
	nor (d438, d333, d354);
	xnor (d439, d382, d385);
	or (d440, d385, d387);
	nand (d441, d335, d344);
	and (d442, d369, d378);
	nand (d443, d358, d364);
	nor (d444, d359, d378);
	nor (d445, d373, d386);
	or (d446, d342, d352);
	or (d447, d350, d382);
	or (d448, d372, d377);
	not (d449, d386);
	xnor (d450, d370, d384);
	nor (d451, d335, d351);
	or (d452, d355, d374);
	not (d453, d165);
	nor (d454, d367, d378);
	or (d455, d343, d386);
	nor (d456, d378, d380);
	nand (d457, d337, d341);
	and (d458, d334, d381);
	xor (d459, d345, d361);
	not (d460, d134);
	or (d461, d345, d386);
	xor (d462, d362, d383);
	buf (d463, d387);
	nor (d464, d352, d387);
	not (d465, d306);
	nand (d466, d340, d384);
	xor (d467, d360, d366);
	and (d468, d336, d345);
	buf (d469, d190);
	nand (d470, d332, d362);
	and (d471, d340, d354);
	not (d472, d225);
	not (d473, d450);
	nand (d474, d399, d442);
	xnor (d475, d400, d402);
	nand (d476, d411, d471);
	and (d477, d396, d437);
	not (d478, d361);
	buf (d479, d196);
	nand (d480, d407, d431);
	not (d481, d370);
	buf (d482, d130);
	nor (d483, d446, d455);
	buf (d484, d363);
	not (d485, d140);
	and (d486, d409, d445);
	xor (d487, d427, d438);
	not (d488, d123);
	and (d489, d438, d445);
	or (d490, d420, d448);
	xor (d491, d427, d462);
	not (d492, d43);
	and (d493, d412, d444);
	buf (d494, d180);
	not (d495, d237);
	nor (d496, d404, d434);
	xnor (d497, d393, d401);
	nand (d498, d401, d460);
	xnor (d499, d448, d456);
	and (d500, d429, d433);
	nand (d501, d426, d435);
	not (d502, d55);
	xnor (d503, d390, d429);
	xor (d504, d440, d464);
	or (d505, d404, d454);
	xor (d506, d429, d463);
	or (d507, d394, d397);
	nand (d508, d389, d455);
	buf (d509, d414);
	buf (d510, x1);
	or (d511, d404, d439);
	not (d512, d126);
	buf (d513, d425);
	nand (d514, d404, d446);
	xnor (d515, d446, d461);
	buf (d516, d369);
	not (d517, d271);
	not (d518, d60);
	assign f1 = d476;
	assign f2 = d478;
	assign f3 = d509;
	assign f4 = d474;
	assign f5 = d483;
	assign f6 = d472;
	assign f7 = d497;
	assign f8 = d510;
	assign f9 = d475;
	assign f10 = d499;
	assign f11 = d517;
	assign f12 = d511;
	assign f13 = d502;
	assign f14 = d514;
	assign f15 = d504;
endmodule
